//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Mon Aug 19 22:28:56 2024

module map_ram (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [4:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [14:0] ada;
input [4:0] din;
input [14:0] adb;

wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [1:1] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [1:1] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [2:2] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [2:2] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [3:3] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [3:3] sdpb_inst_7_dout;
wire [30:0] sdpb_inst_8_dout_w;
wire [4:4] sdpb_inst_8_dout;
wire [30:0] sdpb_inst_9_dout_w;
wire [4:4] sdpb_inst_9_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h00000FFF00000FFF00000FFF00001FFF00001FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h000007FF000007FF000007FF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h000007FF00000FFF00000FFF00001FFF00001FFF00001FFF00001FFF00003FFF;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h000007FF000007FF000007FF000003FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF000007FF;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h000007FF00000FFF00000FFF00000FFF00001FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h000007FF000007FF000007FF000003FF000003FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF000007FF;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h000007FF000007FF00000FFF00000FFF00000FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h000007FF000007FF000007FF000003FF000003FF000003FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h00003FFF00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF000007FF;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h000007FF000007FF000007FF00000FFF00000FFF00000FFF00000FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h000007FF000007FF000007FF000003FF000003FF000003FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h00007FFF00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF000007FF;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h000007FF000007FF000007FF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h000007FF000007FF000007FF000003FF000003FF000003FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h00007FFF00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h000007FF000007FF000007FF000007FF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h000007FF000007FF000007FF000007FF000003FF000003FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h00007FFF00007FFF00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h00000FFF00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h000007FF000007FF000007FF000007FF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h000007FF000007FF000007FF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h00007FFF00007FFF00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h000007FF000007FF000007FF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h00000FFF000007FF000007FF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h00007FFF00007FFF00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF000003FF;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h000007FF000007FF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h00000FFF00000FFF000007FF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h00007FFF00007FFF00007FFF00003FFF00003FFF00001FFF00001FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF000003FF;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000FFFF00007FFF00007FFF00003FFF00003FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000FFFF00007FFF00007FFF00003FFF00003FFF00003FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h00000FFF00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h00000FFF00000FFF00001FFF00001FFF00001FFF00001FFF00001FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000FFFF00007FFF00007FFF00007FFF00003FFF00003FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h00001FFF00000FFF00000FFF00000FFF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000FFFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h00001FFF00001FFF00000FFF00000FFF00000FFF000007FF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000FFFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF000007FF000007FF;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00001FFF;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h00003FFF00003FFF00001FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h00007FFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF00003FFF;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF000007FF;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h00007FFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h00003FFF00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h00007FFF00007FFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h00003FFF00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h00007FFF00007FFF00007FFF00007FFF00007FFF00007FFF00007FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h00003FFF00003FFF00003FFF00007FFF00007FFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h00007FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF00007FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h00003FFF00003FFF00007FFF00007FFF00007FFF00007FFF00007FFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h00003FFF00003FFF00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h00003FFF00003FFF00007FFF00007FFF00007FFF00007FFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h00003FFF00003FFF00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h00003FFF00003FFF00007FFF00007FFF00007FFF0000FFFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h00003FFF00001FFF00001FFF00001FFF00001FFF00001FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h00003FFF00003FFF00007FFF00007FFF00007FFF0000FFFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h00003FFF00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h00003FFF00003FFF00007FFF00007FFF00007FFF0000FFFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00001FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h00003FFF00001FFF00001FFF00001FFF00000FFF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h00003FFF00003FFF00007FFF00007FFF00007FFF0000FFFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00001FFF00001FFF00001FFF;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF000007FF000007FF;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h00001FFF00003FFF00003FFF00007FFF00007FFF0000FFFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00001FFF00001FFF;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h00003FFF00001FFF00001FFF00000FFF00000FFF00000FFF000007FF000007FF;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h00001FFF00003FFF00003FFF00007FFF00007FFF0000FFFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00000FFF00001FFF;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h00001FFF00001FFF00000FFF00000FFF00000FFF000007FF000007FF000007FF;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h0000FFFF0000FFFF0000FFFF0000FFFF00007FFF00007FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h00001FFF00001FFF00003FFF00003FFF00007FFF00007FFF0000FFFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h00000FFF000007FF000007FF000007FF00000FFF00000FFF00000FFF00001FFF;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h00001FFF00001FFF00000FFF00000FFF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h0000FFFF0000FFFF0000FFFF00007FFF00007FFF00007FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h00001FFF00001FFF00003FFF00003FFF00007FFF00007FFF00007FFF0000FFFF;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h000007FF000007FF000007FF000007FF000007FF00000FFF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h00001FFF00001FFF00000FFF00000FFF000007FF000007FF000007FF000007FF;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h0000FFFF0000FFFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h00001FFF00001FFF00001FFF00003FFF00003FFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h000007FF000007FF000007FF000007FF000007FF000007FF00000FFF00000FFF;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h00001FFF00000FFF00000FFF000007FF000007FF000007FF000007FF000003FF;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h00007FFF00007FFF00007FFF00007FFF00007FFF00003FFF00003FFF00001FFF;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h00000FFF00001FFF00001FFF00003FFF00003FFF00007FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h000007FF000007FF000007FF000007FF000007FF000007FF000007FF00000FFF;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h00001FFF00000FFF00000FFF000007FF000007FF000007FF000003FF000003FF;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h00007FFF00007FFF00007FFF00007FFF00003FFF00003FFF00003FFF00001FFF;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h00000FFF00001FFF00001FFF00003FFF00003FFF00003FFF00007FFF00007FFF;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h000007FF000007FF000007FF000007FF000007FF000007FF000007FF00000FFF;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h00003FFC00003FFC00003FFC00007FFC00007FFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h00001FFC00001FFC00001FFC000C1FFC000C1FFC000C1FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h0000FFFC0000FFFC00007FFC00307FFC00003FFC00003FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h00001FFC00003FFC00003FFC00007FFC00007FFC00007FFC00007FFC0000FFFC;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h00001FFC00001FFC000C1FFC000C0FFC000C1FFC000C1FFC000C1FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h0000FFFC0000FFFC00307FFC00307FFC00303FFC00003FFC00003FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h00001FFC00003FFC00003FFC00003FFC00007FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h00001FFC00001FFC00001FFC000C0FFC000C0FFC000C1FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_0B = 256'h0000FFFC0030FFFC00307FFC00307FFC00303FFC00303FFC00003FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_0D = 256'h00001FFC00001FFC00003FFC00003FFC00003FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h00001FFC00001FFC00001FFC00000FFC000C0FFC00000FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h0000FFFC0000FFFC0030FFFC00307FFC00307FFC00003FFC00003FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h00001FFC00001FFC00001FFC00003FFC00003FFC00003FFC00003FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h00001FFC00001FFC00001FFC00000FFC00000FFC00000FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h0001FFFC0000FFFC0000FFFC00307FFC00007FFC00003FFC00003FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h00001FFC00001FFC00001FFC00003FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h00001FFC00001FFC00001FFC00000FFC000C0FFC00000FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_17 = 256'h0001FFFC0000FFFC0000FFFC00007FFC00007FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h00003FFC00003FFC00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_19 = 256'h00001FFC00001FFC00001FFC00001FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h00001FFC00001FFC00001FFC000C1FFC000C0FFC000C0FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h0001FFFC0001FFFC0000FFFC0000FFFC00007FFC00007FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h00003FFC00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h00001FFC00001FFC00001FFC00001FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h00001FFC00001FFC000C1FFC000C1FFC000C1FFC000C1FFC000C1FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h0001FFFC0001FFFC0000FFFC0000FFFC00007FFC00007FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h00001FFC00001FFC00001FFC00003FFC00003FFC00183FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_22 = 256'h00003FFC00001FFC00001FFC000C1FFC000C1FFC000C1FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_23 = 256'h0001FFFC0001FFFC0000FFFC0000FFFC00007FFC00007FFC00003FFC00303FFC;
defparam sdpb_inst_2.INIT_RAM_24 = 256'h00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC00000FFC;
defparam sdpb_inst_2.INIT_RAM_25 = 256'h00001FFC00001FFC00003FFC00003FFC00183FFC00183FFC00183FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_26 = 256'h00303FFC00003FFC00001FFC00001FFC000C1FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_27 = 256'h0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC00007FFC00307FFC00303FFC;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC00000FFC;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h00003FFC00003FFC00003FFC00183FFC00183FFC00183FFC00183FFC00183FFC;
defparam sdpb_inst_2.INIT_RAM_2A = 256'h00303FFC00303FFC00003FFC00001FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h0003FFFC0001FFFC0001FFFC0000FFFC0000FFFC00307FFC00307FFC00307FFC;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h00003FFC00003FFC00003FFC00003FFC00183FFC00183FFC00183FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_2E = 256'h00303FFC00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_2F = 256'h0003FFFC0001FFFC0001FFFC0000FFFC0000FFFC0000FFFC00307FFC00307FFC;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h00003FFC00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h00003FFC00003FFC00007FFC00007FFC00007FFC00187FFC00007FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_32 = 256'h00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h0003FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC00007FFC00307FFC;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h00007FFC00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_35 = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_37 = 256'h0003FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC0000FFFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h00007FFC00007FFC00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h0003FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC0060FFFC0000FFFC;
defparam sdpb_inst_2.INIT_RAM_3C = 256'h00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC00001FFC00001FFC;
defparam sdpb_inst_2.INIT_RAM_3D = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC00007FFC;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h0000FFFC0000FFFC00007FFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h0001FFFC0001FFFC0001FFFC0001FFFC0000FFFC0060FFFC0060FFFC0060FFFC;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h00007FFC00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC00001FFC;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_02 = 256'h0060FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h0001FFFC0001FFFC0001FFFC0001FFFC0060FFFC0060FFFC0060FFFC0060FFFC;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h0000FFFC00007FFC00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_05 = 256'h0001FFFC0001FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_06 = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0001FFFC0001FFFC0001FFFC;
defparam sdpb_inst_3.INIT_RAM_07 = 256'h0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC0060FFFC0060FFFC0060FFFC;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h0000FFFC00007FFC00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_09 = 256'h0001FFFC0001FFFC0001FFFC0001FFFC0001FFFC0001FFFC0001FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_0A = 256'h0000FFFC0000FFFC0000FFFC0001FFFC0001FFFC0001FFFC0001FFFC0001FFFC;
defparam sdpb_inst_3.INIT_RAM_0B = 256'h0001FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0060FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_0C = 256'h0000FFFC0000FFFC00007FFC00007FFC00003FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC0001FFFC0001FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_0E = 256'h0000FFFC0000FFFC0001FFFC0001FFFC0001FFFC0181FFFC0001FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h0000FFFC0000FFFC00007FFC00007FFC00007FFC00003FFC00183FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_11 = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC0001FFFC0001FFFC;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h0000FFFC0000FFFC0001FFFC0001FFFC0181FFFC0181FFFC0183FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_13 = 256'h0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_14 = 256'h0000FFFC0000FFFC00007FFC00007FFC00007FFC00183FFC00183FFC00183FFC;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC00C1FFFC;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h0000FFFC0060FFFC0001FFFC0181FFFC0181FFFC0183FFFC0183FFFC0183FFFC;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h0000FFFC00007FFC00007FFC00007FFC00007FFC00007FFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_18 = 256'h00C0FFFC0000FFFC00007FFC00007FFC00183FFC00183FFC00183FFC00183FFC;
defparam sdpb_inst_3.INIT_RAM_19 = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC00C1FFFC00C1FFFC;
defparam sdpb_inst_3.INIT_RAM_1A = 256'h0060FFFC0060FFFC0061FFFC0001FFFC0181FFFC0183FFFC0183FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_1B = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_1C = 256'h00C0FFFC00C0FFFC00007FFC00187FFC00183FFC00183FFC00183FFC00183FFC;
defparam sdpb_inst_3.INIT_RAM_1D = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0003FFFC00C1FFFC00C1FFFC00C1FFFC;
defparam sdpb_inst_3.INIT_RAM_1E = 256'h0060FFFC0060FFFC0061FFFC0061FFFC0001FFFC0183FFFC0003FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_1F = 256'h00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC00007FFC0060FFFC;
defparam sdpb_inst_3.INIT_RAM_20 = 256'h00C0FFFC00007FFC00007FFC00007FFC00183FFC00183FFC00183FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC00C1FFFC00C0FFFC;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h0060FFFC0060FFFC0061FFFC0001FFFC0001FFFC0003FFFC0003FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_23 = 256'h00003FFC00003FFC00003FFC00003FFC00003FFC00007FFC00007FFC00007FFC;
defparam sdpb_inst_3.INIT_RAM_24 = 256'h0000FFFC00007FFC00007FFC00003FFC00003FFC00183FFC00001FFC00001FFC;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC00C0FFFC;
defparam sdpb_inst_3.INIT_RAM_26 = 256'h00007FFC0060FFFC0000FFFC0001FFFC0001FFFC0003FFFC0003FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC00007FFC00007FFC;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h0000FFFC00007FFC00007FFC00003FFC00003FFC00003FFC00001FFC00001FFC;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC0001FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h00007FFC0000FFFC0000FFFC0001FFFC0001FFFC0003FFFC0003FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC00003FFC00007FFC;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h00007FFC00007FFC00003FFC00003FFC00003FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h0003FFFC0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_2E = 256'h00007FFC00007FFC0000FFFC0000FFFC0001FFFC0001FFFC0003FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h00003FFC00001FFC00001FFC000C1FFC00003FFC00003FFC00003FFC00007FFC;
defparam sdpb_inst_3.INIT_RAM_30 = 256'h00007FFC00007FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_3.INIT_RAM_31 = 256'h0003FFFC0003FFFC0003FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_32 = 256'h00007FFC00007FFC0000FFFC0000FFFC0001FFFC0001FFFC0001FFFC0003FFFC;
defparam sdpb_inst_3.INIT_RAM_33 = 256'h00001FFC00001FFC000C1FFC000C1FFC000C1FFC00003FFC00003FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h00007FFC00007FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h0003FFFC0003FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC0000FFFC;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h00007FFC00007FFC00007FFC0000FFFC0000FFFC0001FFFC0001FFFC0001FFFC;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h00001FFC000C1FFC000C1FFC000C1FFC000C1FFC000C1FFC00003FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_38 = 256'h00007FFC00003FFC00003FFC00001FFC00001FFC00001FFC00001FFC00000FFC;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h0001FFFC0001FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC00007FFC;
defparam sdpb_inst_3.INIT_RAM_3A = 256'h00003FFC00007FFC00007FFC0000FFFC0000FFFC0001FFFC0001FFFC0001FFFC;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h00001FFC00001FFC000C1FFC000C1FFC000C1FFC00001FFC00001FFC00003FFC;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h00007FFC00003FFC00003FFC00001FFC00001FFC00001FFC00000FFC00000FFC;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h0001FFFC0001FFFC0001FFFC0001FFFC0000FFFC0000FFFC0000FFFC00007FFC;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h00003FFC00007FFC00007FFC0000FFFC0000FFFC0000FFFC0001FFFC0001FFFC;
defparam sdpb_inst_3.INIT_RAM_3F = 256'h00001FFC00001FFC00001FFC000C1FFC00001FFC00001FFC00001FFC00003FFC;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_01 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_02 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_03 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_04 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_05 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_06 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_07 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_09 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_0A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_0B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_0C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_0D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_0E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_0F = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_11 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_12 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_13 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_14 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_15 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_16 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_17 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_18 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_19 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_1A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_1B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_1C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_1D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_1E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_1F = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_20 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_21 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_23 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_24 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_25 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_26 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_27 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_28 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_29 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_2A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_2B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_2C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_2D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_2E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_2F = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_30 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_31 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_32 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_33 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_34 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_35 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_36 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_37 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_38 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_39 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_3A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_3B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_3C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_3D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_3E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_4.INIT_RAM_3F = 256'h0000000300000003000000030000000300000003000000030000000300000003;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_01 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_02 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_03 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_04 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_05 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_06 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_07 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_08 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_09 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_0A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_0B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_0C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_0D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_0E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_0F = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_10 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_11 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_12 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_13 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_14 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_15 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_16 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_17 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_18 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_19 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_1A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_1B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_1C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_1D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_1E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_1F = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_20 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_21 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_22 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_23 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_24 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_25 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_26 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_27 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_28 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_29 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_2A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_2B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_2C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_2D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_2E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_2F = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_30 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_31 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_32 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_33 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_34 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_35 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_36 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_37 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_38 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_39 = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_3A = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_3B = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_3C = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_3E = 256'h0000000300000003000000030000000300000003000000030000000300000003;
defparam sdpb_inst_5.INIT_RAM_3F = 256'h0000000300000003000000030000000300000003000000030000000300000003;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_02 = 256'h000000000000000000000000000C0000000C0000000C00000000000000000000;
defparam sdpb_inst_6.INIT_RAM_03 = 256'h0000000000000000000000000030000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_06 = 256'h0000000000000000000C0000000C0000000FE000000C0000000C000000000000;
defparam sdpb_inst_6.INIT_RAM_07 = 256'h0000000000000000003000000030000000300000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0A = 256'h000000000000000000000000000C0000000C0000000C00000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0B = 256'h000000000030000000300000003F800000300000003000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0E = 256'h00000000000000000000000000000000000C0000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0F = 256'h0000000000000000003000000030000000300000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_13 = 256'h0000000000000000000000000030000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_16 = 256'h00000000000000000000000000000000000C0000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1A = 256'h000000000000000000000000000C0000000C0000000C00000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1E = 256'h0000000000000000000C0000000C0000000FE000000C0000000C000000000000;
defparam sdpb_inst_6.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000001800000000000000000000;
defparam sdpb_inst_6.INIT_RAM_22 = 256'h000000000000000000000000000C0000000C0000000C00000000000000000000;
defparam sdpb_inst_6.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000300000;
defparam sdpb_inst_6.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_25 = 256'h0000000000000000000000000000000000180000001800000018000000000000;
defparam sdpb_inst_6.INIT_RAM_26 = 256'h00300000000000000000000000000000000C0000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000030000000300000;
defparam sdpb_inst_6.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_29 = 256'h0000000000000000000000000018000000180000001FC0000018000000180000;
defparam sdpb_inst_6.INIT_RAM_2A = 256'h0030000000300000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2B = 256'h00000000000000000000000000000000000000000030000000300000003F8000;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000180000001800000018000000000000;
defparam sdpb_inst_6.INIT_RAM_2E = 256'h0030000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000030000000300000;
defparam sdpb_inst_6.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000001800000000000000000000;
defparam sdpb_inst_6.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000300000;
defparam sdpb_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000060000000000000;
defparam sdpb_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000006000000060000000600000;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_02 = 256'h0060000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_03 = 256'h000000000000000000000000000000000060000000600000007F000000600000;
defparam sdpb_inst_7.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000006000000060000000600000;
defparam sdpb_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000060000000000000;
defparam sdpb_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000018000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000018000000000000;
defparam sdpb_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_12 = 256'h0000000000000000000000000000000001800000018000000180000000000000;
defparam sdpb_inst_7.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000001800000018000000180000;
defparam sdpb_inst_7.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000C00000;
defparam sdpb_inst_7.INIT_RAM_16 = 256'h000000000060000000000000018000000180000001FC00000180000001800000;
defparam sdpb_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_18 = 256'h00C000000000000000000000000000000018000000180000001FC00000180000;
defparam sdpb_inst_7.INIT_RAM_19 = 256'h00000000000000000000000000000000000000000000000000C0000000C00000;
defparam sdpb_inst_7.INIT_RAM_1A = 256'h0060000000600000006000000000000001800000018000000180000000000000;
defparam sdpb_inst_7.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1C = 256'h00C0000000C00000000000000018000000180000001FC0000018000000180000;
defparam sdpb_inst_7.INIT_RAM_1D = 256'h000000000000000000000000000000000000000000C0000000C0000000FE0000;
defparam sdpb_inst_7.INIT_RAM_1E = 256'h00600000007F0000006000000060000000000000018000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000600000;
defparam sdpb_inst_7.INIT_RAM_20 = 256'h00C0000000000000000000000000000000180000001800000018000000000000;
defparam sdpb_inst_7.INIT_RAM_21 = 256'h00000000000000000000000000000000000000000000000000C0000000C00000;
defparam sdpb_inst_7.INIT_RAM_22 = 256'h0060000000600000006000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000001800000000000000000000;
defparam sdpb_inst_7.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000C00000;
defparam sdpb_inst_7.INIT_RAM_26 = 256'h0000000000600000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2F = 256'h000000000000000000000000000C000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_33 = 256'h0000000000000000000C0000000C0000000C0000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_37 = 256'h00000000000C0000000C0000000FE000000C0000000C00000000000000000000;
defparam sdpb_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3B = 256'h0000000000000000000C0000000C0000000C0000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3F = 256'h000000000000000000000000000C000000000000000000000000000000000000;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[30:0],sdpb_inst_8_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 1;
defparam sdpb_inst_8.BIT_WIDTH_1 = 1;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_8.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[30:0],sdpb_inst_9_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_9.READ_MODE = 1'b0;
defparam sdpb_inst_9.BIT_WIDTH_0 = 1;
defparam sdpb_inst_9.BIT_WIDTH_1 = 1;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_9.RESET_MODE = "SYNC";
defparam sdpb_inst_9.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_9.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(sdpb_inst_2_dout[1]),
  .I1(sdpb_inst_3_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(sdpb_inst_4_dout[2]),
  .I1(sdpb_inst_5_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(sdpb_inst_6_dout[3]),
  .I1(sdpb_inst_7_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_4 (
  .O(dout[4]),
  .I0(sdpb_inst_8_dout[4]),
  .I1(sdpb_inst_9_dout[4]),
  .S0(dff_q_0)
);
endmodule //map_ram
