//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Wed Sep 24 21:24:33 2025

module texture_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [27:0] prom_inst_0_dout_w;
wire [3:0] prom_inst_0_dout;
wire [27:0] prom_inst_1_dout_w;
wire [7:4] prom_inst_1_dout;
wire [27:0] prom_inst_2_dout_w;
wire [11:8] prom_inst_2_dout;
wire [27:0] prom_inst_3_dout_w;
wire [15:12] prom_inst_3_dout;
wire [15:0] prom_inst_4_dout_w;
wire [15:0] prom_inst_4_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[12])
);
defparam lut_inst_0.INIT = 4'h2;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[10]),
  .I2(ad[11]),
  .I3(ad[12])
);
defparam lut_inst_1.INIT = 16'h0200;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],prom_inst_0_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hA66666AA2A0AAA2AAA2AAA626660660A6AA02226222222AAA6666A2022A6666A;
defparam prom_inst_0.INIT_RAM_01 = 256'hAA66660666666AAA0222AAAA226ACA22A066AA0A666AAA66022222666666622A;
defparam prom_inst_0.INIT_RAM_02 = 256'h022AAA22AAA6AAA0AAA22260622662AAA2666AA0A666666A2222222AAA62022A;
defparam prom_inst_0.INIT_RAM_03 = 256'hAA666AAAA2206666A66A22AA66666AAA22AA60666AA0262AA66666226666666A;
defparam prom_inst_0.INIT_RAM_04 = 256'hFEEEEEFF1FDFFF1FFF1FFFE1EEEDEEDFEFFD111EEE1111FFFEEEEF1D11FEEEEF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFEEEEDEEEEEEFFFD111FFFF11EF0F11FDEEFFDFEEEFFFEED11111EEEEEEE11F;
defparam prom_inst_0.INIT_RAM_06 = 256'hD11FFF11FFFEFFFDFFF111EDE11EE1FFF1EEEFFDFEEEEEEF1111111FFFE1D11F;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFEEEFFFF11DEEEEFEEF11FFEEEEEFFF11FFEDEEEF11111FFEEEEE11EEEEEEEF;
defparam prom_inst_0.INIT_RAM_08 = 256'h6555A7649589BA5658674A7C89554969A77766B5866498864A5996645666446D;
defparam prom_inst_0.INIT_RAM_09 = 256'h75A69771454AA85767673C765749435755AA576758735885BA7A79BA79529988;
defparam prom_inst_0.INIT_RAM_0A = 256'h8644998857FC875655457869777675556764446AD44B74688B6546768C777855;
defparam prom_inst_0.INIT_RAM_0B = 256'h559BA88665557A9657CBA96765559988A5C5A9885556AA878554356954467456;
defparam prom_inst_0.INIT_RAM_0C = 256'h75575856555855D55655CCA958577D5B87869CC6775AAB898467789A86877999;
defparam prom_inst_0.INIT_RAM_0D = 256'h997799597799BB779797BB7BB770777BB7775775559799577597D5557795B979;
defparam prom_inst_0.INIT_RAM_0E = 256'h5795799D97B9977970995BB59B7BB79797BB7777755775977577799757979779;
defparam prom_inst_0.INIT_RAM_0F = 256'h5799779970799B79997797BB5757B57999B75B5799787797BB7777777B997957;
defparam prom_inst_0.INIT_RAM_10 = 256'h79B79799B7597BD97B55777B777B577B559B79B750977597B7B7757799B7799B;
defparam prom_inst_0.INIT_RAM_11 = 256'h997799597799BB779797BB7BB770777BB7775775559799577597D7597795B979;
defparam prom_inst_0.INIT_RAM_12 = 256'h5795799D97B9977970995BB59B7BB79797BB7777755775977577799757979779;
defparam prom_inst_0.INIT_RAM_13 = 256'h5799779970799B79997797BB5757B57999B75B5799787797BB7777777B997957;
defparam prom_inst_0.INIT_RAM_14 = 256'hACC4BAF10FAEF3CC02CCA0FF25AFFF4CFF4CC11605C055C164DBACF45EF56CCF;
defparam prom_inst_0.INIT_RAM_15 = 256'hCBAECB041A99AEEFBB211FCCCFF03B0ED0F1F37DAC545EF5DCFF35AAFDAAAA53;
defparam prom_inst_0.INIT_RAM_16 = 256'hF205CCAE054CBACA055CAFFBDCCAF1BA55C9FD55ECA1F0FCCC13D25525B0555C;
defparam prom_inst_0.INIT_RAM_17 = 256'h0C54DAFF4CAF0EA0CAADCFBBBFFEF41CAF1FCF0ECACD0144B005CC5514FB233C;
defparam prom_inst_0.INIT_RAM_18 = 256'h77666677777776669CCCBCC7BB9999CC9CB9B99999BB7BCC9CCCCCC9BCC9999C;
defparam prom_inst_0.INIT_RAM_19 = 256'h7766667776666677CCCCC7999CCCBCCC9999BBBB9CBBB799CBBB799C9CC9999C;
defparam prom_inst_0.INIT_RAM_1A = 256'h76667777766677679BBBBB9999CCBBBC999C7999BBC999999CCCBBBCC97CCCCC;
defparam prom_inst_0.INIT_RAM_1B = 256'h7664677767667777CCCCB9CC9CC999CCB9999BBC9CCCC79BCCCB99799C9CCCCC;
defparam prom_inst_0.INIT_RAM_1C = 256'h3B9CBCBCCCCCBAB66BA9999A998999B35BCBBBAABBBBBAB66667366333666366;
defparam prom_inst_0.INIT_RAM_1D = 256'h7B9CA9CBBC9BD9B33B9BB9CCCC9BC9B36B9BB999AA9BC9B36B9CBBBBBBBBC9B4;
defparam prom_inst_0.INIT_RAM_1E = 256'h5BACBBBBBBBBC9B36B9CB999999BB9A66B9CB9CCCC9BC9B66B9CB9CBBC9BCBB6;
defparam prom_inst_0.INIT_RAM_1F = 256'h63336666636663766BBBBABBAABBBBB43BAAA999999A98B33B9CCCCCCCBCC9B3;
defparam prom_inst_0.INIT_RAM_20 = 256'h7493963963774546947476396396455384749639649337539676766648639664;
defparam prom_inst_0.INIT_RAM_21 = 256'h7376473949396396737257383659647664738636666966567393964766776646;
defparam prom_inst_0.INIT_RAM_22 = 256'h939639539497637384964A535386647474864836648664967366384646487396;
defparam prom_inst_0.INIT_RAM_23 = 256'h7566266646653765637539683476496339863656747665649456395363966393;
defparam prom_inst_0.INIT_RAM_24 = 256'h350159350150000056026B53045A0100A0A6609A00A0370050A0000F000B3502;
defparam prom_inst_0.INIT_RAM_25 = 256'hC0A0A75025B64064BBA00C00440BA02A00B0A03A0B190060120100130A400440;
defparam prom_inst_0.INIT_RAM_26 = 256'h5A00503500006505003B00550B90000B025A020A0301B091A370022022A23017;
defparam prom_inst_0.INIT_RAM_27 = 256'h5A100A55A0300004B2602AC0000BB00C055920A001402B024902201006503601;
defparam prom_inst_0.INIT_RAM_28 = 256'h0355432E42424331822365433333386554343B572221653431A4434432353451;
defparam prom_inst_0.INIT_RAM_29 = 256'h5954233475233533445396332340325F032203634452E2411603522265662624;
defparam prom_inst_0.INIT_RAM_2A = 256'hF22283343334245232D3256743615D545353633322433530344330A356255654;
defparam prom_inst_0.INIT_RAM_2B = 256'h13344273614A034352253F4143342345353445757222E15432552331F4246246;
defparam prom_inst_0.INIT_RAM_2C = 256'h2444323243333334544542322232343455534333223344445434434423443345;
defparam prom_inst_0.INIT_RAM_2D = 256'h4443444422332434444334346323344334333334653223323444333244332323;
defparam prom_inst_0.INIT_RAM_2E = 256'h3344323324334443256413333453333234454234234432223455433444434423;
defparam prom_inst_0.INIT_RAM_2F = 256'h4443534334433445445443332344434443443333334453453432222123444444;
defparam prom_inst_0.INIT_RAM_30 = 256'h77667D67778F6681F120EFF00100013056634333234444456776667667556666;
defparam prom_inst_0.INIT_RAM_31 = 256'h7F0207660178668EF53550EE661F1114F54335E4645F3334436435E3454F3340;
defparam prom_inst_0.INIT_RAM_32 = 256'h774E7EE3EED05777EEE504363303FFFE5F56D35556E355537F67153576F44547;
defparam prom_inst_0.INIT_RAM_33 = 256'h7E660E345F004167D4D055F6E6641502456E334E5344F3766761568E66761576;
defparam prom_inst_0.INIT_RAM_34 = 256'hFEEEEEF67FDFFF1FFF67FFE1EEE6EEDFEFFD111E111111FFFEEEEF1D11FEEEEF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFEEEEDEEEEEEFFFD11166FF66678F11FDEE78DFE78FFFEED11111EEEEEEE11F;
defparam prom_inst_0.INIT_RAM_36 = 256'hD1167F11FFFEFFFDFFF111EDE116E1FFF1EEE6667EEEEEEF11111178FFE1D67F;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFEEEFFFF11DEEEEFEEF11FFEEEEEFFF11FFE66EEFF67E1FFE666787EEEEEEEF;
defparam prom_inst_0.INIT_RAM_38 = 256'h2322234410123331221233111122341132214111222343222211001221111222;
defparam prom_inst_0.INIT_RAM_39 = 256'h1112332212223211122332122134221012335223224211112234233351112121;
defparam prom_inst_0.INIT_RAM_3A = 256'h0122334211121121112345110131111000111100131112110001211221122321;
defparam prom_inst_0.INIT_RAM_3B = 256'h1211100111111322221121221112322121122223222342111112234342132112;
defparam prom_inst_0.INIT_RAM_3C = 256'hFEEEEEFE2FDFFF1FFF02FFE1EEE0EEDFEFFD111E111111FFFEEEEF1D11FEEEEF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFEEEEDEEEEEEFFFD111E0FFE0025F11FDEE25DFE25FFFEED11111EEEEEEE11F;
defparam prom_inst_0.INIT_RAM_3E = 256'hD11E2F11FFFEFFFDFFF111EDE110E1FFF1EEEEEE2EEEEEEF11111125FFE1D02F;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFEEEFFFF11DEEEEFEEF11FFEEEEEFFF11FFEEEEEFFE2E1FFEE00252EEEEEEEF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],prom_inst_1_dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hA88888AABA2AAABAAABAAA8B8882882A8AA2BBB8BBBBBBAAA8888AB2BBA8888A;
defparam prom_inst_1.INIT_RAM_01 = 256'hAA88882888888AAA2BBBAAAABB8A0ABBA288AA2A888AAA882BBBBB8888888BBA;
defparam prom_inst_1.INIT_RAM_02 = 256'h2BBAAABBAAA8AAA2AAABBB828BB88BAAAB888AA2A888888ABBBBBBBAAA8B2BBA;
defparam prom_inst_1.INIT_RAM_03 = 256'hAA888AAAABB28888A88ABBAA88888AAABBAA82888AA2B8BAA88888BB8888888A;
defparam prom_inst_1.INIT_RAM_04 = 256'hEAAAAAEE7E4EEE7EEE7EEEA7AAA4AA4EAEE4777AAA7777EEEAAAAE7477EAAAAE;
defparam prom_inst_1.INIT_RAM_05 = 256'hEEAAAA4AAAAAAEEE4777EEEE77AE1E77E4AAEE4EAAAEEEAA477777AAAAAAA77E;
defparam prom_inst_1.INIT_RAM_06 = 256'h477EEE77EEEAEEE4EEE777A4A77AA7EEE7AAAEE4EAAAAAAE7777777EEEA7477E;
defparam prom_inst_1.INIT_RAM_07 = 256'hEEAAAEEEE774AAAAEAAE77EEAAAAAEEE77EEA4AAAE77777EEAAAAA77AAAAAAAE;
defparam prom_inst_1.INIT_RAM_08 = 256'hE88AAEC48A680AAEA2C04A02266848C6A020EAE84EA6846C4A886AA68EAA44C6;
defparam prom_inst_1.INIT_RAM_09 = 256'hEAACA00A466AA4A0E0CE24EA806642A26A8C8EC08402A42AEA0CE8EA268E8646;
defparam prom_inst_1.INIT_RAM_0A = 256'h4C646664A0E4608A8A6604E8022CEA86EEC644CA646004E20EE86CEE420222A8;
defparam prom_inst_1.INIT_RAM_0B = 256'h688EC44AC6A80A8A820EA6C0EAAA6666A62AA84288ACA82048A40AA8664E266E;
defparam prom_inst_1.INIT_RAM_0C = 256'hAEEAE6EEEEE8EE6EE0AE20EAE8E424EE42608E0E04E88C6A680424AE6E6228AA;
defparam prom_inst_1.INIT_RAM_0D = 256'h66AA66E6AA6622AA6A6A22A22AA3AAA22AAAEAAEEE6A66EAAE6A6EEEAA6E26A6;
defparam prom_inst_1.INIT_RAM_0E = 256'hEA6EA6666A266AA6A366E22E62A22A6A6A22AAAAAEEAAE6AAEAAA66AEA6A6AA6;
defparam prom_inst_1.INIT_RAM_0F = 256'hEA66AA66A3A662A666AA6A22EAEA2EA6662AE2EA66ACAA6A22AAAAAAA266A6EA;
defparam prom_inst_1.INIT_RAM_10 = 256'hA62A6A662AE6A266A2EEAAA2AAA2EAA2EE62A62AE36AAE6A2A2AAEAA662AA662;
defparam prom_inst_1.INIT_RAM_11 = 256'h66AA66E6AA6622AA6A6A22A22AA3AAA22AAAEAAEEE6A66EAAE6A6AE6AA6E26A6;
defparam prom_inst_1.INIT_RAM_12 = 256'hEA6EA6666A266AA6A366E22E62A22A6A6A22AAAAAEEAAE6AAEAAA66AEA6A6AA6;
defparam prom_inst_1.INIT_RAM_13 = 256'hEA66AA66A3A662A666AA6A22EAEA2EA6662AE2EA66ACAA6A22AAAAAAA266A6EA;
defparam prom_inst_1.INIT_RAM_14 = 256'h8003CAE71EA8ED001B02A3EE958EEC10EE10077935237505936C82E158E5902E;
defparam prom_inst_1.INIT_RAM_15 = 256'h2E880E135A66AAACCE957E000EC1FE3A43E7EFF4A07178E760EED5A8E4AAAA5D;
defparam prom_inst_1.INIT_RAM_16 = 256'hE93700881710CA0A15508EEC4008E5C85506E6558287E3E0027D6955B7E15550;
defparam prom_inst_1.INIT_RAM_17 = 256'h105148EE12AE3AA32AA60EEEEEEAE172AE5C0E3A28043731C335005571ECBDF0;
defparam prom_inst_1.INIT_RAM_18 = 256'hEEAAAAEEEEEEEAAA2CCC8CCE882222CC2C8282222288E8CC2CCCCCC28CC2222C;
defparam prom_inst_1.INIT_RAM_19 = 256'hEEAAAAEEEAAAAAEECCCCCE222CCC8CCC222288882C888E22C888E22C2CC2222C;
defparam prom_inst_1.INIT_RAM_1A = 256'hEAAAEEEEEAAAEEAE2888882222CC888C222CE22288C222222CCC888CC2ECCCCC;
defparam prom_inst_1.INIT_RAM_1B = 256'hEAAEAEEEA0AA0EEECCCC82CC2CC222CC8222288C2CCCCE28CCC822E22C2CCCCC;
defparam prom_inst_1.INIT_RAM_1C = 256'h682CACACCCCC848AA822222602E2008668AA88648888868ACAAC6AA6668AA6AA;
defparam prom_inst_1.INIT_RAM_1D = 256'hE82C42A88C282286682A82CCAA08A286A80A82224428C086A82CA88888A8C06E;
defparam prom_inst_1.INIT_RAM_1E = 256'h884CA8886886C266882CA22222288268A80C82CCCCE6C08AAA0C80C88A28C88A;
defparam prom_inst_1.INIT_RAM_1F = 256'hA666AAAAA68AA6CAA88882884488888E6646422E22242E86682ACCCCCA8CC286;
defparam prom_inst_1.INIT_RAM_20 = 256'h0AE8C86C880086CCCE0E086C88C8A646AE0EC88C8AC84C88EA0C0888AAC8CAAC;
defparam prom_inst_1.INIT_RAM_21 = 256'hC808E06CAC8CA8CAC8042068686AAE0888086A8AA88C8A4A06C8CAAC8A008AAA;
defparam prom_inst_1.INIT_RAM_22 = 256'hC6AA8E44CACC8808AACA8E4866A8A80C0AAAAA6AAAAC8CEA08AA68AA8AAAC8CA;
defparam prom_inst_1.INIT_RAM_23 = 256'h08A848AA88A6808488086C888E0A8A866EAA886CCE08A4CAC86A6A88A4CA86C6;
defparam prom_inst_1.INIT_RAM_24 = 256'hD70576D505700000590B9E5F01780700A08B906A00A0DD0350A0000E000CF70B;
defparam prom_inst_1.INIT_RAM_25 = 256'h00808D5097CB30B1EC800200310C80B830C0A0D80E7603905907007D08300110;
defparam prom_inst_1.INIT_RAM_26 = 256'h580350D70000B70700DC00550C40000E097A0B0A0D07C067AFD009B09BABD07D;
defparam prom_inst_1.INIT_RAM_27 = 256'h7A70087580D00001C990B820003EC0020576B08005309C093609B0500970D905;
defparam prom_inst_1.INIT_RAM_28 = 256'hDBFFF974B5D5B9737757FDFBBB99771B1B99BFDF757BDB9B93B9B9BF97BFBBDF;
defparam prom_inst_1.INIT_RAM_29 = 256'hD5BD793BBF5B9D9B7BDBBF9779DDBF9AFB55FB599B17F5D313F5D733FDFF7F7F;
defparam prom_inst_1.INIT_RAM_2A = 256'h8577D9BB9B7BFFD3B9DB71537911D0BD17BB5BBB73999D9DB977BDF79F7BD19D;
defparam prom_inst_1.INIT_RAM_2B = 256'h19BB953B11DFD9F7B5FD9AD1DB59577B5D9FDD5B577563DD75DB59BFAD5D37B1;
defparam prom_inst_1.INIT_RAM_2C = 256'h5BBFB597B9779B9DFDDFF79753359B7B111BD79B33379B9B1F9DB7BB579D97DD;
defparam prom_inst_1.INIT_RAM_2D = 256'h9BB99FBB55795B7B99B79D99F75B7BB79999775B3D7339957BBF99B5DB995B79;
defparam prom_inst_1.INIT_RAM_2E = 256'hB79B75773B77BBD95F1D3BD99BD799B39BBFB77D39DB75759DFFDB999BB99B79;
defparam prom_inst_1.INIT_RAM_2F = 256'hBBD9F9B779B7BBD1BBFBB99557D9D9DDDBB97B779579D7BD9D9535737BD9B9BB;
defparam prom_inst_1.INIT_RAM_30 = 256'h55FF5AF155523F71CF53CC01F311F571FFF799773579997D1551115115DBF11F;
defparam prom_inst_1.INIT_RAM_31 = 256'h3C1315111335F15CCB9DD1EAFD323559CBB99DEB1BD2B779B7FB7DC7DFD27993;
defparam prom_inst_1.INIT_RAM_32 = 256'h33DE1CC9EEA1D333AEED1B9F9937EEECDCDFC7BDBFE9DDD73E155D9911EB9D93;
defparam prom_inst_1.INIT_RAM_33 = 256'h3E3F3C9DDC11B311AB81DD0FAD193D139DFC779CB997E7FFD1F39F3C11313DF1;
defparam prom_inst_1.INIT_RAM_34 = 256'hEAAAAAEAEE4EEE7EEEAEEEA7AAAAAA4EAEE4777A777777EEEAAAAE7477EAAAAE;
defparam prom_inst_1.INIT_RAM_35 = 256'hEEAAAA4AAAAAAEEE4777AAEEAAAE2E77E4AAE24EAE2EEEAA477777AAAAAAA77E;
defparam prom_inst_1.INIT_RAM_36 = 256'h477AEE77EEEAEEE4EEE777A4A77AA7EEE7AAAAAAEAAAAAAE777777E2EEA74AEE;
defparam prom_inst_1.INIT_RAM_37 = 256'hEEAAAEEEE774AAAAEAAE77EEAAAAAEEE77EEAAAAAEEAEA7EEAAAAE2EAAAAAAAE;
defparam prom_inst_1.INIT_RAM_38 = 256'hACAAAC00626ACCC6AA6ACC6666AAC066CAA60666AAAC0CAAAA66226AA6666AAA;
defparam prom_inst_1.INIT_RAM_39 = 256'h666ACCAA6AAACA666AACCA6AA6C0AA626ACC4AACAA0A6666AAC0ACCC4666A6A6;
defparam prom_inst_1.INIT_RAM_3A = 256'h26AACC0A666A66A666AC046626C66662226666226C666A662226A66AA66AACA6;
defparam prom_inst_1.INIT_RAM_3B = 256'h6A66622666666CAAAA66A6AA666ACAA6A66AAAACAAAC0A66666AAC0C0A6CA66A;
defparam prom_inst_1.INIT_RAM_3C = 256'hEAAAAAE67E4EEE7EEED7EEA7AAADAA4EAEE4777A777777EEEAAAAE7477EAAAAE;
defparam prom_inst_1.INIT_RAM_3D = 256'hEEAAAA4AAAAAAEEE47776DEE6DD71E77E4AA714EA71EEEAA477777AAAAAAA77E;
defparam prom_inst_1.INIT_RAM_3E = 256'h47767E77EEEAEEE4EEE777A4A77DA7EEE7AAA6667AAAAAAE77777771EEA74D7E;
defparam prom_inst_1.INIT_RAM_3F = 256'hEEAAAEEEE774AAAAEAAE77EEAAAAAEEE77EEA66AAEE67A7EEA6DD717AAAAAAAE;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],prom_inst_2_dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h2111112242022242224222141110110212204441444444222111124044211112;
defparam prom_inst_2.INIT_RAM_01 = 256'h2211110111111222044422224412324420112202111222110444441111111442;
defparam prom_inst_2.INIT_RAM_02 = 256'h0442224422212220222444101441142224111220211111124444444222140442;
defparam prom_inst_2.INIT_RAM_03 = 256'h2211122224401111211244221111122244221011122041422111114411111112;
defparam prom_inst_2.INIT_RAM_04 = 256'hB33333BBCBBBBBCBBBCBBB3C333B33BB3BBBCCC333CCCCBBB3333BCBCCB3333B;
defparam prom_inst_2.INIT_RAM_05 = 256'hBB3333B333333BBBBCCCBBBBCC3B4BCCBB33BBBB333BBB33BCCCCC3333333CCB;
defparam prom_inst_2.INIT_RAM_06 = 256'hBCCBBBCCBBB3BBBBBBBCCC3B3CC33CBBBC333BBBB333333BCCCCCCCBBB3CBCCB;
defparam prom_inst_2.INIT_RAM_07 = 256'hBB333BBBBCCB3333B33BCCBB33333BBBCCBB3B333BCCCCCBB33333CC3333333B;
defparam prom_inst_2.INIT_RAM_08 = 256'hC44C5C44D45DE5C4C5C5C5DEDD4CCDCD55D5C4DCD4CCD5DCC5CDD4CC44CCCCCE;
defparam prom_inst_2.INIT_RAM_09 = 256'hCCDCD55BC4455D45C5C4CE4C4545C4C544554C454D54C5D4D5DDC555DD43DD5D;
defparam prom_inst_2.INIT_RAM_0A = 256'hDCCCDDDDC566D54C4C44D54DD5D44CC4CCCCCCC5E4CE5C455DC4CC44D655DD4C;
defparam prom_inst_2.INIT_RAM_0B = 256'h4C5DDD5CC4C455DCCD6D5DC544CCDD5554645D5544CC55D554CCCCC544C4D444;
defparam prom_inst_2.INIT_RAM_0C = 256'hA99A9D9C999599B9954966D5959D5E9DD5D5556C5D955DD5D45D5D5DDCD55555;
defparam prom_inst_2.INIT_RAM_0D = 256'h33AA3393AA33CCAA3A3ACCACCAA4AAACCAAA9AA9993A339AA93AB999AA39C3A3;
defparam prom_inst_2.INIT_RAM_0E = 256'h9A39A33B3AC33AA3A4339CC93CACCA3A3ACCAAAAA99AA93AA9AAA33A9A3A3AA3;
defparam prom_inst_2.INIT_RAM_0F = 256'h9A33AA33A4A33CA333AA3ACC9A9AC9A333CA9C9A33A2AA3ACCAAAAAAAC33A39A;
defparam prom_inst_2.INIT_RAM_10 = 256'hA3CA3A33CA93ACB3AC99AAACAAAC9AAC993CA3CA943AA93ACACAA9AA33CAA33C;
defparam prom_inst_2.INIT_RAM_11 = 256'h33AA3393AA33CCAA3A3ACCACCAA4AAACCAAA9AA9993A339AA93ABA93AA39C3A3;
defparam prom_inst_2.INIT_RAM_12 = 256'h9A39A33B3AC33AA3A4339CC93CACCA3A3ACCAAAAA99AA93AA9AAA33A9A3A3AA3;
defparam prom_inst_2.INIT_RAM_13 = 256'h9A33AA33A4A33CA333AA3ACC9A9AC9A333CA9C9A33A2AA3ACCAAAAAAAC33A39A;
defparam prom_inst_2.INIT_RAM_14 = 256'h2335A2BC4B23BC33443324BB4D2BBB53BB533CC54D34DD3C55BA23B5D3BD533B;
defparam prom_inst_2.INIT_RAM_15 = 256'h3A233A45C2AA233BAA4CCB333BB4CA43B4BCBCDB23D5D3BDB3BBCD22BB2222DC;
defparam prom_inst_2.INIT_RAM_16 = 256'hB44D33234D53A2324DD32BBAB332BCA2DD3ABBDD332CB4B333CCB4DD4DA4DDD3;
defparam prom_inst_2.INIT_RAM_17 = 256'h43D5B2BB532B4324322B3BAAABB3B5C32BCB3B43323B4C55A44D33DDC5BA4CC3;
defparam prom_inst_2.INIT_RAM_18 = 256'h22AAAA2222222AAACCCC4CC244CCCCCCCC4C4CCCCC4424CCCCCCCCCC4CCCCCCC;
defparam prom_inst_2.INIT_RAM_19 = 256'h22AAAA222AAAAA22CCCCC2CCCCCC4CCCCCCC4444CC4442CCC4442CCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_1A = 256'h2AAA22222AAA22A2C44444CCCCCC444CCCCC2CCC44CCCCCCCCCC444CCC2CCCCC;
defparam prom_inst_2.INIT_RAM_1B = 256'h2AA9A222ABAAB222CCCC4CCCCCCCCCCC4CCCC44CCCCCC2C4CCC4CC2CCCCCCCCC;
defparam prom_inst_2.INIT_RAM_1C = 256'h94CCCCCCCCCC444AA44CCCC4CC3CCC4924CC444C4444444AAAAA9AA9992AA9AA;
defparam prom_inst_2.INIT_RAM_1D = 256'h24CCC4C44CC4DC4994CC4CCCCCC4CC49A4CC4CCC44C4CC49A4CCC44444C4CC49;
defparam prom_inst_2.INIT_RAM_1E = 256'h244CC4444444CC49A4CCCCCCCCC44C42A4CC4CCCCCB4CC4AACCC4CC44CC4CC4A;
defparam prom_inst_2.INIT_RAM_1F = 256'hA999AAAAA9AAA9AAA4444C44CC44444994444C4BCCC4CB4994CCCCCCCC4CCC49;
defparam prom_inst_2.INIT_RAM_20 = 256'hB1B9BA9BA9BB121AB9B9B29B29BA12A939B9BA9B21B99A29BABAB2A213A9BAA1;
defparam prom_inst_2.INIT_RAM_21 = 256'hA9B29B9B1B9BA9BAA9B1AB939A23A9BA21B9BA9AA2AB2AAAB9B9BA1A2ABB2A1A;
defparam prom_inst_2.INIT_RAM_22 = 256'hB93A9BA9B1BA29B931BA1BA92932A1B1B13A139AA13A21BAB9AA931A1A1329BA;
defparam prom_inst_2.INIT_RAM_23 = 256'hB2A212AA1AA29BAA29B29BA399BA13299B3A922AA9BAAAA1B12A9329A9BA29B9;
defparam prom_inst_2.INIT_RAM_24 = 256'hCD0CDACD0CD00000D5045ADC05D20C00202550A20020CD04D020000B000ACD04;
defparam prom_inst_2.INIT_RAM_25 = 256'h30202DD04DA55055AA200300550A204240A020C20ACA0450C40C00CC02500550;
defparam prom_inst_2.INIT_RAM_26 = 256'hD204D0CD00005D0D00CA00DD0AA0000A04D204020C0CA0AC2CD004404424C0CD;
defparam prom_inst_2.INIT_RAM_27 = 256'hD2C002DD20C00005A4504230004AA0030DDA40200C504A045A0440C005D0C50C;
defparam prom_inst_2.INIT_RAM_28 = 256'hDE6E6E65E6E6EE6EF6EEE66EEE6E6FF6FEEEEF66666D66EEEE7EEEE6E6E6E665;
defparam prom_inst_2.INIT_RAM_29 = 256'h6F6E666EF66EE66EEE6EFE666E6DEDED5E6E5E76EEF6FEEEEF5666E6E6EE6E66;
defparam prom_inst_2.INIT_RAM_2A = 256'hD666FEEEEE6ED66EE6FE6777E6F66D6EF66EFEEE66EEE6E5EEE6E5F6EE666FE6;
defparam prom_inst_2.INIT_RAM_2B = 256'h66EEE67EF6EF56666ED66DEE6E6EE6E66666E67676665E6E66666EE5D66EF6EF;
defparam prom_inst_2.INIT_RAM_2C = 256'h6EE6E6E66EE6EEE666E666666EEEEE6EF77E66EEEEE6E6EEF666E6EE66E6E666;
defparam prom_inst_2.INIT_RAM_2D = 256'hEEEEE6EE666EEE6EEEE6E6EE666E6EE6EEEE6E6EF66EEEE66EE66EE66EE66E6E;
defparam prom_inst_2.INIT_RAM_2E = 256'hE6EE6666E6E6EE6E66F6EEEEEE66E6EEEEE6E666EE6E666666666EEEEE6EEE6E;
defparam prom_inst_2.INIT_RAM_2F = 256'hEEEE66E66E6EEE6FEE6EE6E6E6EE6E666EEE6E66666EE6E6E6E6E66E6EEEEEEE;
defparam prom_inst_2.INIT_RAM_30 = 256'h77667D6F777EF67E55EE55665E6E56666666EE66E66EEE66F77FFF7FF7666FFE;
defparam prom_inst_2.INIT_RAM_31 = 256'hF5EE67FF6EF7EF755E6E665D6EEEEEEE5EEEE65EFE6EE666E66E665E66EE6EEE;
defparam prom_inst_2.INIT_RAM_32 = 256'hFF65F55E55DE6FFF555EEEE6EEE65555E5E656E6EE5E6666F5F766EEFF5EE6EF;
defparam prom_inst_2.INIT_RAM_33 = 256'hF5FEE5E66566EEF7DED66EE6DE7EE66EEE656665EEE65666676EEEF5FFFFE66F;
defparam prom_inst_2.INIT_RAM_34 = 256'hB33333B19BBBBBCBBB19BB3C333133BB3BBBCCC3CCCCCCBBB3333BCBCCB3333B;
defparam prom_inst_2.INIT_RAM_35 = 256'hBB3333B333333BBBBCCC11BB11192BCCBB3392BB392BBB33BCCCCC3333333CCB;
defparam prom_inst_2.INIT_RAM_36 = 256'hBCC19BCCBBB3BBBBBBBCCC3B3CC13CBBBC3331119333333BCCCCCC92BB3CB19B;
defparam prom_inst_2.INIT_RAM_37 = 256'hBB333BBBBCCB3333B33BCCBB33333BBBCCBB31133BB193CBB31119293333333B;
defparam prom_inst_2.INIT_RAM_38 = 256'h0800081180808888008088888800818880081888000818000088008008888000;
defparam prom_inst_2.INIT_RAM_39 = 256'h8880880080008088800880800881008080889008001088880081088898880808;
defparam prom_inst_2.INIT_RAM_3A = 256'h0800881088808808880819880888888000888800888880880008088008800808;
defparam prom_inst_2.INIT_RAM_3B = 256'h8088800888888800008808008880800808800008000810888880081810880880;
defparam prom_inst_2.INIT_RAM_3C = 256'hB33333BCDBBBBBCBBBCDBB3C333C33BB3BBBCCC3CCCCCCBBB3333BCBCCB3333B;
defparam prom_inst_2.INIT_RAM_3D = 256'hBB3333B333333BBBBCCCCCBBCCCD6BCCBB33D6BB3D6BBB33BCCCCC3333333CCB;
defparam prom_inst_2.INIT_RAM_3E = 256'hBCCCDBCCBBB3BBBBBBBCCC3B3CCC3CBBBC333CCCD333333BCCCCCCD6BB3CBCDB;
defparam prom_inst_2.INIT_RAM_3F = 256'hBB333BBBBCCB3333B33BCCBB33333BBBCCBB3CC33BBCD3CBB3CCCD6D3333333B;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[27:0],prom_inst_3_dout[15:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 4;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h5333335595055595559555393330330535509993999999555333359099533335;
defparam prom_inst_3.INIT_RAM_01 = 256'h5533330333333555099955559935659950335505333555330999993333333995;
defparam prom_inst_3.INIT_RAM_02 = 256'h0995559955535550555999303993395559333550533333359999999555390995;
defparam prom_inst_3.INIT_RAM_03 = 256'h5533355559903333533599553333355599553033355093955333339933333335;
defparam prom_inst_3.INIT_RAM_04 = 256'h7777777787677787778777787776776777768887778888777777778688777777;
defparam prom_inst_3.INIT_RAM_05 = 256'h7777776777777777688877778877878876777767777777776888887777777887;
defparam prom_inst_3.INIT_RAM_06 = 256'h6887778877777776777888767887787778777776777777778888888777786887;
defparam prom_inst_3.INIT_RAM_07 = 256'h7777777778867777777788777777777788777677778888877777778877777777;
defparam prom_inst_3.INIT_RAM_08 = 256'h5555866575778856575648686755475786665685665477654857765456554459;
defparam prom_inst_3.INIT_RAM_09 = 256'h6575766345588656565649655657445655885666566457658868688867547776;
defparam prom_inst_3.INIT_RAM_0A = 256'h6544776656A96655555567676666655556544458954864677855456679666655;
defparam prom_inst_3.INIT_RAM_0B = 256'h5488877555556875569887566555777785958777555588667554455855466556;
defparam prom_inst_3.INIT_RAM_0C = 256'h7557565555575565565599775756695866667995665888676566667765666777;
defparam prom_inst_3.INIT_RAM_0D = 256'h997799597799BB779797BB7BB778777BB777577555979957759765557795B979;
defparam prom_inst_3.INIT_RAM_0E = 256'h5795799697B9977978995BB59B7BB79797BB7777755775977577799757979779;
defparam prom_inst_3.INIT_RAM_0F = 256'h5799779978799B79997797BB5757B57999B75B5799777797BB7777777B997957;
defparam prom_inst_3.INIT_RAM_10 = 256'h79B79799B7597B697B55777B777B577B559B79B758977597B7B7757799B7799B;
defparam prom_inst_3.INIT_RAM_11 = 256'h997799597799BB779797BB7BB778777BB777577555979957759767597795B979;
defparam prom_inst_3.INIT_RAM_12 = 256'h5795799697B9977978995BB59B7BB79797BB7777755775977577799757979779;
defparam prom_inst_3.INIT_RAM_13 = 256'h5799779978799B79997797BB5757B57999B75B5799777797BB7777777B997957;
defparam prom_inst_3.INIT_RAM_14 = 256'h566A557887577966896658779A5777A677A6688B8A68AA68BA65567AA77AB667;
defparam prom_inst_3.INIT_RAM_15 = 256'h6557658A854457775598876667789587687879B656AAA77A66779A55765555A9;
defparam prom_inst_3.INIT_RAM_16 = 256'h798A66578AA655658AA6577566657855AA6476AA76587876668969AA9A58AAA6;
defparam prom_inst_3.INIT_RAM_17 = 256'h86AA6577A65787586556675557777A8657876787656688AA588A66AA8A759996;
defparam prom_inst_3.INIT_RAM_18 = 256'h77666677777776669BBBBBB7BB9999BB9BB9B99999BB7BBB9BBBBBB9BBB9999B;
defparam prom_inst_3.INIT_RAM_19 = 256'h7766667776666677BBBBB7999BBBBBBB9999BBBB9BBBB799BBBB799B9BB9999B;
defparam prom_inst_3.INIT_RAM_1A = 256'h76667777766677679BBBBB9999BBBBBB999B7999BBB999999BBBBBBBB97BBBBB;
defparam prom_inst_3.INIT_RAM_1B = 256'h7664677767667777BBBBB9BB9BB999BBB9999BBB9BBBB79BBBBB99799B9BBBBB;
defparam prom_inst_3.INIT_RAM_1C = 256'h3B9BBBBBBBBBBAB66BA9999A999999B36BBBBBBABBBBBBB66666366333666366;
defparam prom_inst_3.INIT_RAM_1D = 256'h7B9BAABBBB9BC9B33B9BB9BBBB9BB9B36B9BB999AA9BB9B36B9BBBBBBBBBB9B4;
defparam prom_inst_3.INIT_RAM_1E = 256'h6BABBBBBBBBBB9B36B9BB999999BB9B66B9BB9BBBB9BB9B66B9BB9BBBB9BBAB6;
defparam prom_inst_3.INIT_RAM_1F = 256'h63336666636663666BBBBABBAABBBBB43BAAA9A9999A99B33B9BBBBBBBBBB9B3;
defparam prom_inst_3.INIT_RAM_20 = 256'h7493963963774646947476396396465394749639649336639676766649639664;
defparam prom_inst_3.INIT_RAM_21 = 256'h6376473949396396637357393669647664738636666966567393964666776646;
defparam prom_inst_3.INIT_RAM_22 = 256'h9396395394966373949649536396647474964936649664967366394646497396;
defparam prom_inst_3.INIT_RAM_23 = 256'h7666366646663765637639693476496339963666647665649466396363966393;
defparam prom_inst_3.INIT_RAM_24 = 256'h9A08A49A08A00000AB09B5A90AA50800505BB04500509B08A050000700059A09;
defparam prom_inst_3.INIT_RAM_25 = 256'h60505BA09A5BA0BA55500600AA05509580505095058408B08908008905A00AA0;
defparam prom_inst_3.INIT_RAM_26 = 256'hA508A09A0000BA0A009500AA0540000509A509050908504859B009909959908B;
defparam prom_inst_3.INIT_RAM_27 = 256'hA58005AA5090000A59B09560008550060AA4905008A09509A40990800BA09B08;
defparam prom_inst_3.INIT_RAM_28 = 256'hBDEEEDDBDDDDDDDCFDCDEEEDDDDDDFEEEDDDDFEEDDDBEEDDDCFDDDDEDDDEDEEC;
defparam prom_inst_3.INIT_RAM_29 = 256'hEEEDDDDDFEDDDEDDDDEDFEDDDDEBDCDBCDDCCDFDDDEDFCDCCECDEDCDEEEEDEDE;
defparam prom_inst_3.INIT_RAM_2A = 256'hBDDDFDDDDDDDCEECDDFDDEFFDDECEAEDEDEDEDDDDDDDDEDCDDDDDCFDDEDEEEDE;
defparam prom_inst_3.INIT_RAM_2B = 256'hCDDDDDFDECDFCDEDECCEDBDCEDDDCDDEDEDEDEFEFDDDBCEDDDEEDDDCBEDDEDDE;
defparam prom_inst_3.INIT_RAM_2C = 256'hDDDEDDDDEDDDDDDEEEDEEDDDDCCCDDDDEEEDEDDDCCCDDEDDEEDEDDDDDDDEDDEE;
defparam prom_inst_3.INIT_RAM_2D = 256'hDDDDDEDDDDDDCDDDDDDDDEDDEDDDDDDDDDDDDDDDEEDCCDDDDDDEDDDDEDDDDDDD;
defparam prom_inst_3.INIT_RAM_2E = 256'hDDDDDDDDCEDDDDEDDEEECDDDDDEDDDDCDDDEDDDECDEDDDDDDEEEEDDDDDEDDDDD;
defparam prom_inst_3.INIT_RAM_2F = 256'hDDDDEDDDDDEDDDEEDDEDDDDDCDDDEDEEEDDDDDDDDDDDDDDEDEDDCDDCDDDDDDDD;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFEEFBEEFFFCEEFCCCCCCCCCCCCCCDDCEEEDDDDDCDDDDDDEEFFEEEFEEFEEEEEE;
defparam prom_inst_3.INIT_RAM_31 = 256'hECCCCFEECCEFEEFCCDDDECCBEDCCCCCDCDDDDECDEDECDDDDDDEDDECDEEDCDDDC;
defparam prom_inst_3.INIT_RAM_32 = 256'hEEECECCDCCBCEEEECCCDCDDEDDCDCCCCDCDECDDEDECDEEEDECEFDEDDEECDDEDE;
defparam prom_inst_3.INIT_RAM_33 = 256'hECEECCDEECCCDCEEBDBCEDCEBDEDCECCDDECDDDCDDDDCDEEEEECDEECEEEECEEE;
defparam prom_inst_3.INIT_RAM_34 = 256'h7777777337677787773377787773776777768887888888777777778688777777;
defparam prom_inst_3.INIT_RAM_35 = 256'h7777776777777777688833773333478876773467734777776888887777777887;
defparam prom_inst_3.INIT_RAM_36 = 256'h6883378877777776777888767883787778777333377777778888883477786337;
defparam prom_inst_3.INIT_RAM_37 = 256'h7777777778867777777788777777777788777337777337877733334377777777;
defparam prom_inst_3.INIT_RAM_38 = 256'h1111112200011110110111000011120011102000111121111100000110000111;
defparam prom_inst_3.INIT_RAM_39 = 256'h0001111101111100011111011012110001112111112100001112111120001010;
defparam prom_inst_3.INIT_RAM_3A = 256'h0011112100010010001122000010000000000000010001000000100110011110;
defparam prom_inst_3.INIT_RAM_3B = 256'h0100000000000111110010110001111010011111111121000001112121011001;
defparam prom_inst_3.INIT_RAM_3C = 256'h7777777AD767778777BD7778777B776777768887888888777777778688777777;
defparam prom_inst_3.INIT_RAM_3D = 256'h77777767777777776888AB77ABBDE7887677DE677DE777776888887777777887;
defparam prom_inst_3.INIT_RAM_3E = 256'h688AD7887777777677788876788B787778777AAAD7777777888888DE77786BD7;
defparam prom_inst_3.INIT_RAM_3F = 256'h7777777778867777777788777777777788777AA7777AD78777ABBDED77777777;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[15:0],prom_inst_4_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 16;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hBDD7BDD7BDD7BDD7BDD7C638C618C618C618C638C618BDF7BDD7B5B6B5B6BDF7;
defparam prom_inst_4.INIT_RAM_01 = 256'hBDF7E73CE73CE73CE73CE73CE73CE73CEF7DEF7DEF7DEF7DEF5DEF5DEF5DCE59;
defparam prom_inst_4.INIT_RAM_02 = 256'hBDF7E73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CC638;
defparam prom_inst_4.INIT_RAM_03 = 256'hB596D6BAD6BADEDBDEDBE71CE71CE71CE71CDEFBDEFBDEFBDEFBDEFBDEFBB5B6;
defparam prom_inst_4.INIT_RAM_04 = 256'hBDF7E73CE73CE73CE73CE73CE73CEF7DEF7DEF7DF79EEF7DEF7DEF7DF79EC638;
defparam prom_inst_4.INIT_RAM_05 = 256'hBDF7E73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CC638;
defparam prom_inst_4.INIT_RAM_06 = 256'hB596DEDBDEDBDEDBDEDBDEDBE71CE71CE71CE71CDEDBDEFBDEFBDEFBDEFBBDD7;
defparam prom_inst_4.INIT_RAM_07 = 256'hBDF7E73CE73CE73CE73CE73CE73CE73CEF5DEF5DEF5DEF5DEF7DEF7DF79EC638;
defparam prom_inst_4.INIT_RAM_08 = 256'hBDF7E73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CC638;
defparam prom_inst_4.INIT_RAM_09 = 256'hB596DEFBD6BAD6BADEDBDEDBE71CDEFBDEFBE71CE71CE71CDEFBDEFBDEFBB5B6;
defparam prom_inst_4.INIT_RAM_0A = 256'hBDF7E73CE73CE73CE73CEF7DEF7DEF7DEF7DF79EF79EF79EF79EF79EF79EC638;
defparam prom_inst_4.INIT_RAM_0B = 256'hBDD7E73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CC638;
defparam prom_inst_4.INIT_RAM_0C = 256'hB596DEDBD6BADEDBDEDBDEDBE71CE71CE71CE71CDEFBDEFBDEFBDEFBDEFBB5B6;
defparam prom_inst_4.INIT_RAM_0D = 256'hBDD7E73CE73CE73CE73CE73CE73CEF7DF79EF79EF79EF79EEF7DF79EF79EC638;
defparam prom_inst_4.INIT_RAM_0E = 256'hBDD7E73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CE73CC638;
defparam prom_inst_4.INIT_RAM_0F = 256'hB5B6B5B6B5B6B5B6BDF7BDF7BDF7BDF7B5B6BDD7BDD7BDD7BDD7BDD7BDD7BDF7;
defparam prom_inst_4.INIT_RAM_10 = 256'h18A118A118A118A1084018A118A1084008400840188118A118A1084018A118A1;
defparam prom_inst_4.INIT_RAM_11 = 256'h1881B48BBCAC2922AB88AB88AB88AB68AB88AB88AB88AB882902B46AB48B18A1;
defparam prom_inst_4.INIT_RAM_12 = 256'h18A1B48B2102A347A347A347A347A388A347A3479B27A347A34720E2B48B0840;
defparam prom_inst_4.INIT_RAM_13 = 256'h08402902A34751C451A451C44943496351C451C451C4496351A4A368290218A1;
defparam prom_inst_4.INIT_RAM_14 = 256'h18A1AB88A34751C4B3A99AC64943AB88AB8851A4A2E69AC651C4A347AB881061;
defparam prom_inst_4.INIT_RAM_15 = 256'h18A1AB88A34751A49AC68A854983A34792A54122A347AB8851C4A347AB880840;
defparam prom_inst_4.INIT_RAM_16 = 256'h0840AB88A34751A44943498351C4496351A451A4498351A451A4A347AB880840;
defparam prom_inst_4.INIT_RAM_17 = 256'h18A1AB88A34751C4AB68A36751A4AB88AB8851C4A347AB8859C4A347AB880840;
defparam prom_inst_4.INIT_RAM_18 = 256'h18A1B3A9A34751C4AB88A34751C4AB88AB8851A4A347AB8851C49AC6AB8818A1;
defparam prom_inst_4.INIT_RAM_19 = 256'h18A1AB88A34751C451A4498351C4496351C451C4498351A449638A65B3A918A1;
defparam prom_inst_4.INIT_RAM_1A = 256'h18A1AB88A34751C4B3A9A34741228A85A3474983A3479AC64943A347AB881881;
defparam prom_inst_4.INIT_RAM_1B = 256'h1881AB88A36851C4B3A99AC651A4AB88AB8851A4B3889AC651C4A347AB880840;
defparam prom_inst_4.INIT_RAM_1C = 256'h08402902A34751A451C451C451C451C451C451A4494351C451C4A34729020840;
defparam prom_inst_4.INIT_RAM_1D = 256'h0840B46B2102A388A368A347A3479B47A347A347A347A368A34720E2B48B0840;
defparam prom_inst_4.INIT_RAM_1E = 256'h18A1B48BB48B2902AB88AB68AB88AB88AB68AB68B3A9AB882902B48BB48B1061;
defparam prom_inst_4.INIT_RAM_1F = 256'h18A108400840084018A151225122512251224902512218A118A1084018A118A1;
defparam prom_inst_4.INIT_RAM_20 = 256'h18A1BCCCBCCCBCCCBCCC2922B3A959635963B3A929229C299C299C299C2918A1;
defparam prom_inst_4.INIT_RAM_21 = 256'h18A1BCCCB48B9C29B48B9C292102596359632102B48BB48B72E7B48BBCCC18A1;
defparam prom_inst_4.INIT_RAM_22 = 256'h18A1BCCCBCCC72E7B48BBCCCBCCC29222902B48B9C297AC69C299C29BCCC18A1;
defparam prom_inst_4.INIT_RAM_23 = 256'h18A172E728E128E128E141A472E718A118A172E772E749E449E46AA66AA618A1;
defparam prom_inst_4.INIT_RAM_24 = 256'h18A172C728E172C728E17AC69C2929222102BCCCBCCC9C297AC69C299C2918A1;
defparam prom_inst_4.INIT_RAM_25 = 256'h18A1628628E128E128E19B47B48B29022102BCCCB48BB48B28E172E79C2918A1;
defparam prom_inst_4.INIT_RAM_26 = 256'h18A172E7B5B6DEDBDEDB49E49C2921022102BCCCBCCCBCCC28E1BCCCBCCC18A1;
defparam prom_inst_4.INIT_RAM_27 = 256'h18A141C4B5B6DEDBFFFF6AA672E718A118A16AA66AA66AA628E16AA672E718A1;
defparam prom_inst_4.INIT_RAM_28 = 256'h18A172E7B5B6DEDB72C7B48BB48B292229229C2972E7B5B628E1BCCCBCCC18A1;
defparam prom_inst_4.INIT_RAM_29 = 256'h18A16286B5B6FFFF72E79C299C2921022902B48B72E7B5B6DEDBB5B69C2918A1;
defparam prom_inst_4.INIT_RAM_2A = 256'h18A172C7B5B6DEDBB48BB48B9C29210218A19C2972E7B5B672C772C7B48B18A1;
defparam prom_inst_4.INIT_RAM_2B = 256'h18A141A3B5B6290272E772E772E718A110616AA641A341A372E772E76AA618A1;
defparam prom_inst_4.INIT_RAM_2C = 256'h18A172E7FFFF9B479C299C299C29210218A1BCCC9C29BCCCA387BCCCBCCC18A1;
defparam prom_inst_4.INIT_RAM_2D = 256'h18A1628662869C299C29B48BB48B29222102BCCCBCCCBCCCA38772E79C2918A1;
defparam prom_inst_4.INIT_RAM_2E = 256'h18A1BCCCBCCCBCCCB48B9C29BCCC29222102BCCCBCCC9C297AC69C29BCCC18A1;
defparam prom_inst_4.INIT_RAM_2F = 256'h18A16AA66AA649E46AA672E772E718A118A17B076AA66AA67B0772E772E718A1;
defparam prom_inst_4.INIT_RAM_30 = 256'h18A1BCCCBCCCBCCCBCCC2922B3A959635963B3A929229C299C299C299C2918A1;
defparam prom_inst_4.INIT_RAM_31 = 256'h18A1BCCCB48B9C29B48B9C292102596359632102B48BB48B72E7B48BBCCC18A1;
defparam prom_inst_4.INIT_RAM_32 = 256'h18A1BCCCBCCC72E7B48BBCCCBCCC29222902B48B9C297AC69C299C29BCCC18A1;
defparam prom_inst_4.INIT_RAM_33 = 256'h18A172E76AA66AA66AA641A472E718A118A172E772E749E449E46AA66AA618A1;
defparam prom_inst_4.INIT_RAM_34 = 256'h18A1B48BB48BB48B72E77AC69C2929222102BCCCBCCC9C297AC69C299C2918A1;
defparam prom_inst_4.INIT_RAM_35 = 256'h18A19C299C299C29B48B9B47B48B29022102BCCC28E1B48B28E172E79C2918A1;
defparam prom_inst_4.INIT_RAM_36 = 256'h18A1BCCCBCCCBCCCBCCC49E49C292102210272E728E172E728E1BCCCBCCC18A1;
defparam prom_inst_4.INIT_RAM_37 = 256'h18A172E76AA66AA641A46AA672E718A118A16AA66AA6DEDB6AA66AA672E718A1;
defparam prom_inst_4.INIT_RAM_38 = 256'h18A1BCCCBCCCBCCCB48BB48BB48B292229226286DEDB72E7DEDBBCCCBCCC18A1;
defparam prom_inst_4.INIT_RAM_39 = 256'h18A19C299C29BCCC72E79C299C292102290272C7B5B66286B5B69C299C2918A1;
defparam prom_inst_4.INIT_RAM_3A = 256'h18A1B48BB48B9B47B48BB48B9C29210218A19C29BCCCBCCCB48BB48BB48B18A1;
defparam prom_inst_4.INIT_RAM_3B = 256'h18A16AA66AA641A472E772E772E718A110616AA66AA66AA672E772E76AA618A1;
defparam prom_inst_4.INIT_RAM_3C = 256'h18A1BCCC72E79B479C299C299C29210218A1BCCC9C29BCCCA387BCCCBCCC18A1;
defparam prom_inst_4.INIT_RAM_3D = 256'h18A19C299C299C299C29B48BB48B29222102BCCCBCCCBCCCA38772E79C2918A1;
defparam prom_inst_4.INIT_RAM_3E = 256'h18A1BCCCBCCCBCCCB48B9C29BCCC29222102BCCCBCCC9C297AC69C29BCCC18A1;
defparam prom_inst_4.INIT_RAM_3F = 256'h18A16AA66AA649E46AA672E772E718A118A17B076AA66AA67B0772E772E718A1;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_4 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_4_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(dout[1]),
  .I0(prom_inst_0_dout[1]),
  .I1(prom_inst_4_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[2]),
  .I0(prom_inst_0_dout[2]),
  .I1(prom_inst_4_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_19 (
  .O(dout[3]),
  .I0(prom_inst_0_dout[3]),
  .I1(prom_inst_4_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_24 (
  .O(dout[4]),
  .I0(prom_inst_1_dout[4]),
  .I1(prom_inst_4_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[5]),
  .I0(prom_inst_1_dout[5]),
  .I1(prom_inst_4_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_34 (
  .O(dout[6]),
  .I0(prom_inst_1_dout[6]),
  .I1(prom_inst_4_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_39 (
  .O(dout[7]),
  .I0(prom_inst_1_dout[7]),
  .I1(prom_inst_4_dout[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(dout[8]),
  .I0(prom_inst_2_dout[8]),
  .I1(prom_inst_4_dout[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_49 (
  .O(dout[9]),
  .I0(prom_inst_2_dout[9]),
  .I1(prom_inst_4_dout[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_54 (
  .O(dout[10]),
  .I0(prom_inst_2_dout[10]),
  .I1(prom_inst_4_dout[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_59 (
  .O(dout[11]),
  .I0(prom_inst_2_dout[11]),
  .I1(prom_inst_4_dout[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_64 (
  .O(dout[12]),
  .I0(prom_inst_3_dout[12]),
  .I1(prom_inst_4_dout[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_69 (
  .O(dout[13]),
  .I0(prom_inst_3_dout[13]),
  .I1(prom_inst_4_dout[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_74 (
  .O(dout[14]),
  .I0(prom_inst_3_dout[14]),
  .I1(prom_inst_4_dout[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_79 (
  .O(dout[15]),
  .I0(prom_inst_3_dout[15]),
  .I1(prom_inst_4_dout[15]),
  .S0(dff_q_0)
);
endmodule //texture_rom
