module ram_char (
	input  [6:0]   raddr,
	output [511:0] rdata
);

reg [511:0] ram[127:0];
assign rdata = ram[raddr];

initial
begin
	ram[0] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[1] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[2] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[3] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[4] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[5] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[6] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[7] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[8] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[9] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[10] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[11] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[12] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[13] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[14] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[15] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[16] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[17] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[18] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[19] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[20] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[21] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[22] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[23] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[24] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[25] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[26] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[27] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[28] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[29] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[30] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[31] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[32] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[33] = 512'h00000000000000000000000003C003C003C003C003C003C001C001800180018001800180018001800180000000000000018003C003C001800000000000000000;
	ram[34] = 512'h000000000318073807380E700C6018C0318021000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[35] = 512'h000000000000000000000000040804080408040804087FFE7FFE7FFE0810081008100810081008107FFE7FFE7FFE183010201020102010200000000000000000;
	ram[36] = 512'h00000000000000000100010003C00D3009181918193819381D000D000F00070003C001E001F00130013801183918391831183130196007C00100010001000000;
	ram[37] = 512'h00000000000000000000000038106C104420C620C640C640C640C680C68044806D38396C024402C602C604C604C608C608C60844106C10380000000000000000;
	ram[38] = 512'h0000000000000000000000000F0019003180318031803180310033003A001C00387C3C104C10CE10C620C720C320C1C0C1C260E6317C1E380000000000000000;
	ram[39] = 512'h0000000038003C003C000C000C000800300060000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[40] = 512'h000000000002000400080018003000200060004000C000C001800180018001800180018001800180018000C000C0004000600020003000180008000400020000;
	ram[41] = 512'h0000000040002000100018000C0004000600020003000300018001800180018001800180018001800180030003000300060004000C0018001000200040000000;
	ram[42] = 512'h0000000000000000000000000000000000C001C001C030C6388E1C9C06B001C001C006B01C9C388E318601C001C001C000000000000000000000000000000000;
	ram[43] = 512'h00000000000000000000000000000000000000800080008000800080008000803FFE008000800080008000800080008000000000000000000000000000000000;
	ram[44] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038003C003C000C000C00080030006000;
	ram[45] = 512'h00000000000000000000000000000000000000000000000000000000000000007FFE000000000000000000000000000000000000000000000000000000000000;
	ram[46] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018003C003C0018000000000000000000;
	ram[47] = 512'h000000000000000200060004000C000800180010003000200060004000C000800180010003000200060004000C00080018001000300020006000400000000000;
	ram[48] = 512'h00000000000000000000000003C006200C30181818181808300C300C300C300C300C300C300C300C300C300C1808181818180C30062003C00000000000000000;
	ram[49] = 512'h000000000000000000000000008001801F800180018001800180018001800180018001800180018001800180018001800180018003C01FF80000000000000000;
	ram[50] = 512'h00000000000000000000000007E008381018200C200C300C300C000C001800180030006000C0018003000200040408041004200C3FF83FF80000000000000000;
	ram[51] = 512'h00000000000000000000000007C018603030301830183018001800180030006003C0007000180008000C000C300C300C30083018183007C00000000000000000;
	ram[52] = 512'h0000000000000000000000000060006000E000E0016001600260046004600860086010603060206040607FFC0060006000600060006003FC0000000000000000;
	ram[53] = 512'h0000000000000000000000000FFC0FFC10001000100010001000100013E0143018181008000C000C000C000C300C300C20182018183007C00000000000000000;
	ram[54] = 512'h00000000000000000000000001E006180C180818180010001000300033E0363038183808300C300C300C300C300C180C18080C180E3003E00000000000000000;
	ram[55] = 512'h0000000000000000000000001FFC1FFC100830102010202000200040004000400080008001000100010001000300030003000300030003000000000000000000;
	ram[56] = 512'h00000000000000000000000007E00C301818300C300C300C380C38081E180F2007C018F030783038601C600C600C600C600C3018183007C00000000000000000;
	ram[57] = 512'h00000000000000000000000007C01820301030186008600C600C600C600C600C701C302C186C0F8C000C0018001800103030306030C00F800000000000000000;
	ram[58] = 512'h0000000000000000000000000000000000000000000000000000018003C003C001800000000000000000000000000000018003C003C001800000000000000000;
	ram[59] = 512'h00000000000000000000000000000000000000000000000000000000038003800380000000000000000000000000000000000380038003800180030003000000;
	ram[60] = 512'h00000000000000000000000000040008001000200040008001000200040008001000100008000400020001000080004000200010000800040000000000000000;
	ram[61] = 512'h00000000000000000000000000000000000000000000000000007FFE000000000000000000007FFE000000000000000000000000000000000000000000000000;
	ram[62] = 512'h00000000000000000000000020001000080004000200010000800040002000100008000800100020004000800100020004000800100020000000000000000000;
	ram[63] = 512'h00000000000000000000000003E00C18180C10063006380638063806000C0018007000C0008000800080008000000000018003C003C001800000000000000000;
	ram[64] = 512'h00000000000000000000000003E006100C08180430D431B221326332632266226622662266626664666426E8333030021004180C0C1803E00000000000000000;
	ram[65] = 512'h000000000000000000000000038003800380038004C004C004C004C00C4008600860086018201FF0103010301030201820182018601CF83E0000000000000000;
	ram[66] = 512'h0000000000000000000000007FE018381818180C180C180C180C180C181818301FE01818180C180418061806180618061806180C18187FF00000000000000000;
	ram[67] = 512'h00000000000000000000000003E0061C080C180630023002300060006000600060006000600060006000600030023002100418080C1003E00000000000000000;
	ram[68] = 512'h0000000000000000000000007FC0187018181808180C180C1806180618061806180618061806180618061804180C180C1818181818607FC00000000000000000;
	ram[69] = 512'h0000000000000000000000007FFC180C180418021802180018001810181018301FF0183018101810180018001800180218021804180C7FFC0000000000000000;
	ram[70] = 512'h0000000000000000000000007FFC181C180418021802180018001810181018301FF018301810181018101800180018001800180018007E000000000000000000;
	ram[71] = 512'h00000000000000000000000003C00C300810181830083008200060006000600060006000607E60186018201830183018101818180C2007C00000000000000000;
	ram[72] = 512'h000000000000000000000000FC3F300C300C300C300C300C300C300C300C300C3FFC300C300C300C300C300C300C300C300C300C300CFC3F0000000000000000;
	ram[73] = 512'h0000000000000000000000001FF8018001800180018001800180018001800180018001800180018001800180018001800180018001801FF80000000000000000;
	ram[74] = 512'h00000000000000000000000007FE006000600060006000600060006000600060006000600060006000600060006000600060006000600060706070C071803F00;
	ram[75] = 512'h0000000000000000000000007E7C183018201860184018801880190019001B001D801D8018C018C018601860183018301830181818187E3E0000000000000000;
	ram[76] = 512'h0000000000000000000000007E001800180018001800180018001800180018001800180018001800180018001800180218021804180C7FFC0000000000000000;
	ram[77] = 512'h000000000000000000000000F00F381C381C381C381C382C2C2C2C2C2C2C2C4C2C4C264C264C264C268C228C238C238C230C230C210CF13F0000000000000000;
	ram[78] = 512'h000000000000000000000000F01F380438042C042C0426042604230423042184218420C420C42064206420342034201C201C200C200CF8040000000000000000;
	ram[79] = 512'h00000000000000000000000003C00C3018181008300C300C6004600660066006600660066006600660062006300C300C100818180C3003C00000000000000000;
	ram[80] = 512'h0000000000000000000000007FF01818180C180618061806180618061806180C18181FE01800180018001800180018001800180018007E000000000000000000;
	ram[81] = 512'h00000000000000000000000003C00C3018181008300C300C6006600660066006600660066006600660066006278438CC386C18780C7003E00032003C001C0000;
	ram[82] = 512'h0000000000000000000000007FE018381818180C180C180C180C180C181818301FE018C018C0186018601860183018301830181818187E1E0000000000000000;
	ram[83] = 512'h0000000000000000000000000FC818783018601860086008600070003C001F0007C001F000780018001C400C400C600C200C3018383027E00000000000000000;
	ram[84] = 512'h0000000000000000000000003FFC3184218641824182018001800180018001800180018001800180018001800180018001800180018007E00000000000000000;
	ram[85] = 512'h000000000000000000000000FC3E30083008300830083008300830083008300830083008300830083008300830083008300818101C2007C00000000000000000;
	ram[86] = 512'h0000000000000000000000007C1E180C1808180818080C100C100C100C100C200620062006200640034003400340038001800180010001000000000000000000;
	ram[87] = 512'h000000000000000000000000F3CF618661842184208430C431C431C431C831C811C812481A681A681A701C700C700C700C300C20082008200000000000000000;
	ram[88] = 512'h0000000000000000000000007C3E180818100C100C20062006400340038001800180018001C002C0026004600470083008301818101C7C3E0000000000000000;
	ram[89] = 512'h0000000000000000000000007E3E3808180818100C100C100C200620062003400340038001800180018001800180018001800180018007E00000000000000000;
	ram[90] = 512'h0000000000000000000000001FFE1C0C180C3018201800300060006000C000C00180018003000300060006000C00180218063004301C7FFC0000000000000000;
	ram[91] = 512'h00000000000003FC030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003FC00000000;
	ram[92] = 512'h000000000000000000001800180008000C0004000600060002000300010001800180008000C000400060006000300030003000180018000C000C000C00060000;
	ram[93] = 512'h0000000000003FC000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C000C03FC000000000;
	ram[94] = 512'h0000000003C003E00620081000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[95] = 512'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFF;
	ram[96] = 512'h000000001E0003000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[97] = 512'h000000000000000000000000000000000000000000000000000007E01830301830183018003807D81C183018601860186018601930791F8E0000000000000000;
	ram[98] = 512'h000000000000000000000800780018001800180018001800180019E01A381C181C0C180C180C180C180C180C180C180C18081C181C3013E00000000000000000;
	ram[99] = 512'h000000000000000000000000000000000000000000000000000003E00E100C1818183018300030003000300030003004180418080C1003E00000000000000000;
	ram[100] = 512'h000000000000000000000008007800180018001800180018001807D80C38181818183018301830183018301830183018101818380C5E07900000000000000000;
	ram[101] = 512'h000000000000000000000000000000000000000000000000000003C00C3008181808300C300C300C3FFC300030003000180418080E1803E00000000000000000;
	ram[102] = 512'h000000000000000000000000007C0186010603060300030003003FF803000300030003000300030003000300030003000300030003001FF00000000000000000;
	ram[103] = 512'h000000000000000000000000000000000000000000000000000003EE0C36081818181818181808180C300FE0180018001FC00FF8181C300C300C300C181807E0;
	ram[104] = 512'h000000000000000000000800780018001800180018001800180019E01A301C18181818181818181818181818181818181818181818187E7E0000000000000000;
	ram[105] = 512'h000000000000000000000000018003C0018000000000000000801F8001800180018001800180018001800180018001800180018001801FF80000000000000000;
	ram[106] = 512'h000000000000000000000000003800780030000000000000001003F0003000300030003000300030003000300030003000300030003000300030186018400F80;
	ram[107] = 512'h0000000000000000000008007800180018001800180018001800187C183018201840188019801B801EC01CC01860183018301818181C7E3E0000000000000000;
	ram[108] = 512'h0000000000000000000000801F80018001800180018001800180018001800180018001800180018001800180018001800180018001801FF80000000000000000;
	ram[109] = 512'h0000000000000000000000000000000000000000000000002000EF3C71C6618661866186618661866186618661866186618661866186F3CF0000000000000000;
	ram[110] = 512'h000000000000000000000000000000000000000000000000000009E07A301C18181818181818181818181818181818181818181818187E7E0000000000000000;
	ram[111] = 512'h000000000000000000000000000000000000000000000000000003C00C3008181818100C300C300C300C300C300C300C181818180C3003C00000000000000000;
	ram[112] = 512'h000000000000000000000000000000000000000000000000000009E07A301C181808180C180C180C180C180C180C180C18181C181E3019E01800180018007E00;
	ram[113] = 512'h000000000000000000000000000000000000000000000000000003C80C78183818183018301830183018301830183018101818380C780798001800180018007E;
	ram[114] = 512'h0000000000000000000000801F80018001800180018001800180018001800180018001800180018001800180018001800180018001801FF80000000000000000;
	ram[115] = 512'h000000000000000000000000000000000000000000000000000003E4061C0C0C0C040C040E0007C001F00078001C100C100C180C1C1813F00000000000000000;
	ram[116] = 512'h00000000000000000000000000000000010001000100030007003FF8030003000300030003000300030003000300030003040304018800F00000000000000000;
	ram[117] = 512'h000000000000000000000000000000000000000000000000080878781818181818181818181818181818181818181818181818380C5E07900000000000000000;
	ram[118] = 512'h00000000000000000000000000000000000000000000000000007C3E180C180818180C100C100420062006200340034003C00180018001000000000000000000;
	ram[119] = 512'h0000000000000000000000000000000000000000000000000000FBCF618621843184318431C811C81AC81A481A700E700C700C300C2004200000000000000000;
	ram[120] = 512'h00000000000000000000000000000000000000000000000000003E7C0C100E100620034003400180018001C0026004600430081818187C7E0000000000000000;
	ram[121] = 512'h00000000000000000000000000000000000000000000000000007C3E1818181008100C100420062006200240034001400180018001000100010002003E003C00;
	ram[122] = 512'h00000000000000000000000000000000000000000000000000003FF830383030206020E000C001800380030006000E040C04180C30183FF80000000000000000;
	ram[123] = 512'h00000000000C00100020002000200020002000200020002000200020002000C001800040002000200020002000200020002000200020002000200010000C0000;
	ram[124] = 512'h00800080008000800080008000800080008000800080008000800080008000800080008000800080008000800080008000800080008000800080008000800080;
	ram[125] = 512'h000000001800040002000200020002000200020002000200020002000200018000C0010002000200020002000200020002000200020002000200040018000000;
	ram[126] = 512'h00001E0023004182408200E400380000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ram[127] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end

endmodule

