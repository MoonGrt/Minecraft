//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Mon Apr 01 19:39:52 2024

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [23:0] dout;
input clk;
input oce;
input ce;
input reset;
input [7:0] ad;

wire [7:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[7:0],dout[23:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[7:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 32;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000BFB50000C2B80000BCB20000ADA00000ADA00000ADA00000ADA00000ADA0;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000BDB3001ECFC70019CEC6000ACAC20000C7BE0000C4BA0000BCB20000BDB3;
defparam prom_inst_0.INIT_RAM_02 = 256'h0082E4E00082E4E00087E5E10082E4E0006EE0DB0064DED90064DED90000BDB3;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000BFB50073E1DC0078E2DE007DE3DF0082E4E00082E4E0007DE3DF007DE3DF;
defparam prom_inst_0.INIT_RAM_04 = 256'h008CE7E3008CE7E3008CE7E30091E8E4008CE7E3008CE7E3008CE7E30000C3B9;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000BFB5005ADCD60069DFDA0078E2DE0087E5E1008CE7E30087E5E10087E5E1;
defparam prom_inst_0.INIT_RAM_06 = 256'h0096E9E5009BEAE60091E8E4008CE7E3008CE7E30091E8E40091E8E40000C5BC;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000BFB5007DE3DF007DE3DF007DE3DF0082E4E00082E4E00087E5E10091E8E4;
defparam prom_inst_0.INIT_RAM_08 = 256'h0091E8E40091E8E40096E9E50087E5E10091E8E4008CE7E30096E9E50000C4BA;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000C3B90073E1DC0073E1DC0078E2DE007DE3DF0082E4E00091E8E40091E8E4;
defparam prom_inst_0.INIT_RAM_0A = 256'h0087E5E10082E4E00082E4E00069DFDA0069DFDA0091E8E4009BEAE60000C4BA;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000C3B9007DE3DF007DE3DF0087E5E10087E5E10087E5E10087E5E10087E5E1;
defparam prom_inst_0.INIT_RAM_0C = 256'h0082E4E00082E4E00073E1DC0082E4E00082E4E00087E5E10091E8E40000C4BA;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000C1B7006EE0DB007DE3DF0087E5E10087E5E10082E4E00087E5E10087E5E1;
defparam prom_inst_0.INIT_RAM_0E = 256'h0069DFDA0069DFDA0069DFDA0069DFDA0082E4E0008CE7E3009BEAE60000C4BA;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000BFB5005FDDD70073E1DC0082E4E0007DE3DF0073E1DC006EE0DB0069DFDA;
defparam prom_inst_0.INIT_RAM_10 = 256'h0069DFDA0069DFDA0069DFDA00A0EBE80082E4E000A0EBE80096E9E50000C5BC;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000BBB0003CD5CF0055DBD50069DFDA0069DFDA0069DFDA0069DFDA0069DFDA;
defparam prom_inst_0.INIT_RAM_12 = 256'h0096E9E50091E8E40096E9E50096E9E50082E4E000A5ECE90096E9E50000C6BD;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000C1B70082E4E0008CE7E30096E9E5009BEAE6009BEAE60096E9E50096E9E5;
defparam prom_inst_0.INIT_RAM_14 = 256'h00A5ECE900A5ECE900A0EBE800A5ECE900AAEDEA00AAEDEA00A5ECE90000C6BD;
defparam prom_inst_0.INIT_RAM_15 = 256'h0000B8AD0064DED90087E5E1009BEAE600A0EBE8009BEAE600A0EBE800A0EBE8;
defparam prom_inst_0.INIT_RAM_16 = 256'h00A5ECE900AAEDEA00AAEDEA00AAEDEA00AAEDEA00AAEDEA00AAEDEA0000C7BE;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000B2A60023D0C8003CD5CF005FDDD70087E5E1009BEAE6009BEAE600A0EBE8;
defparam prom_inst_0.INIT_RAM_18 = 256'h00A0EBE800AAEDEA00AAEDEA00A5ECE900A0EBE800A0EBE800AAEDEA0000C7BE;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000B2A60000C8BF0005C9C10019CEC60050DAD40078E2DE008CE7E30096E9E5;
defparam prom_inst_0.INIT_RAM_1A = 256'h009BEAE600A0EBE800A0EBE800A0EBE80091E8E40096E9E500A5ECE90000C7BE;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000B1A5000FCBC3000FCBC3001ECFC7002DD2CB0046D7D10078E2DE008CE7E3;
defparam prom_inst_0.INIT_RAM_1C = 256'h007DE3DF0082E4E00087E5E10082E4E0007DE3DF008CE7E30096E9E50000C6BD;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000AC9F0000C1B70000C2B80000C5BC000FCBC30032D3CC006EE0DB0078E2DE;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000C1B70000C7BE0000C1B70000C1B70000C1B70000C1B70000C1B70000C1B7;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000BBB00000BEB40000C2B80000C5BC0000C6BD0000C6BD0005C9C10000C2B8;

endmodule //Gowin_pROM
