//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.02
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Thu Aug 29 10:35:20 2024

module texture_rom (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire [27:0] prom_inst_2_dout_w;
wire [27:0] prom_inst_3_dout_w;
wire [27:0] prom_inst_4_dout_w;
wire [27:0] prom_inst_5_dout_w;
wire [27:0] prom_inst_6_dout_w;
wire [27:0] prom_inst_7_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFF0FFFFF0FF00000FF0FFFFF0FFF0F00F0FFF0FF00F0FF0FF0F0000F000FFF0F;
defparam prom_inst_0.INIT_RAM_25 = 256'hF0F0FFF0FFFFF0FFFFF00F00FF0FF0FFF0F0F0FF0FFF0FF0FF0F00FF0FF00FF0;
defparam prom_inst_0.INIT_RAM_26 = 256'hFF0FF0FF0000FF0F00FF00FF0FF0000F0FFF0F0F0F0FF0FFFFF00FF0FFFFF0FF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFF00FFFF0F0000FFFF0FFF000FFF00F0FFFF0F00FF0FF0FFF0FF0F00FF0FF0F;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_24 = 256'hFF0FFFFF0FF00000FF0FFFFF0FFF0F00F0FFF0FF00F0FF0FF0F0000F000FFF0F;
defparam prom_inst_1.INIT_RAM_25 = 256'hF0F0FFF0FFFFF0FFFFF00F00FF0FF0FFF0F0F0FF0FFF0FF0FF0F00FF0FF00FF0;
defparam prom_inst_1.INIT_RAM_26 = 256'hFF0FF0FF0000FF0F00FF00FF0FF0000F0FFF0F0F0F0FF0FFFFF00FF0FFFFF0FF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFF00FFFF0F0000FFFF0FFF000FFF00F0FFFF0F00FF0FF0FFF0FF0F00FF0FF0F;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hF44444FFFF8FFFFFFFFFFF4F4448448F4FF8FFF444FFFFFFF4444FF8FFF4444F;
defparam prom_inst_2.INIT_RAM_01 = 256'hFF44448444444FFF8FFFFFFFFF4F0FFFF844FF8F444FFF448FFFFF4444444FFF;
defparam prom_inst_2.INIT_RAM_02 = 256'h8FFFFFFFFFF4FFF8FFFFFF484FF44FFFFF444FF8F444444FFFFFFFFFFF4F8FFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hFF444FFFFFF84444F44FFFFF44444FFFFFFF48444FFFFFFFF44444FF4444444F;
defparam prom_inst_2.INIT_RAM_04 = 256'h5C9E3945BE7CC3F5F11922C019AC1D2C3BE951AF1615B64323EDB4079700311B;
defparam prom_inst_2.INIT_RAM_05 = 256'hBF01E9BF196111DB6948F790CA692DFD8E04C969C09CF40DB3E6CF83F997DA74;
defparam prom_inst_2.INIT_RAM_06 = 256'h2253A952FA8659A0BF68D46ECDF39FD868054312C45CB462097C538772BCE1DD;
defparam prom_inst_2.INIT_RAM_07 = 256'h88E9766018C982E0CF0C4A3B7DFEBC67382D2E4299D0301B3CF1CF0F9626B786;
defparam prom_inst_2.INIT_RAM_08 = 256'hAACAAAAACA9AACCAAC99AAACAAAC9AAC99ACAACA97AAA9AACACAA9AAAACAAAAC;
defparam prom_inst_2.INIT_RAM_09 = 256'hAAAAAA9AAAAACCAAAAAACCACCAA7AAACCAAA9AA999AAAA9AA9AACA9AAAA9CAAA;
defparam prom_inst_2.INIT_RAM_0A = 256'h9AA9AAACAACAAAAAA7AA9CC9ACACCAAAAACCAAAAA99AA9AAA9AAAAAA9AAAAAAA;
defparam prom_inst_2.INIT_RAM_0B = 256'h9AAAAAAAA7AAACAAAAAAAACC9A9AC9AAAACA9C9AAAA4AAAACCAAAAAAACAAAA9A;
defparam prom_inst_2.INIT_RAM_0C = 256'h322586FF1F61DB22372465FF292FFA02FF332ED06977C92906DA24E290F9024D;
defparam prom_inst_2.INIT_RAM_0D = 256'h7D323D1796CD6479AE18DF222EA2CE7787FFFEF862D2E2CFF2FFA950F8666699;
defparam prom_inst_2.INIT_RAM_0E = 256'hF15F22132E22A61629910FFA9220F9B2992EFC99260DF7F225CBC0996CD19992;
defparam prom_inst_2.INIT_RAM_0F = 256'h129390FF376F7746566C2FCFDEF4F2C66F8A2D4460187E62A449229BF3D979E2;
defparam prom_inst_2.INIT_RAM_10 = 256'h7333337777777777777777373337337737777773777777777333377777733337;
defparam prom_inst_2.INIT_RAM_11 = 256'h7733337333333777777777777737377777337777333777337777773333333777;
defparam prom_inst_2.INIT_RAM_12 = 256'h7777777777737777777777373773377777333777733333377777777777377777;
defparam prom_inst_2.INIT_RAM_13 = 256'h7733377777773333733777773333377777773733377773777333337733333337;
defparam prom_inst_2.INIT_RAM_14 = 256'h77111177777771113DDD5DD555AAAADD3D5A5AAAAA5555DD3DDDDDDA5DDAAAAD;
defparam prom_inst_2.INIT_RAM_15 = 256'h7711117771111177DDDDD5AA3DDD5DDDAAAA55553D5555AAD5555AAD3DDAAAAD;
defparam prom_inst_2.INIT_RAM_16 = 256'h7111777771117717355555AAAADD555D3AAD5AAA55DAAAAA3DDD555DDA5DDDDD;
defparam prom_inst_2.INIT_RAM_17 = 256'h711E177719119777DDDD5ADD3DDAAADD5AAAA55D3DDDD5A5DDD5AA5A3DADDDDD;
defparam prom_inst_2.INIT_RAM_18 = 256'h9933339999999333D222A229AADDDD22D2ADADDDDDAA9A22D222222DA22DDDD2;
defparam prom_inst_2.INIT_RAM_19 = 256'h9933339993333399222229DDD222A222DDDDAAAAD2AAA9DD2AAA9DD2D22DDDD2;
defparam prom_inst_2.INIT_RAM_1A = 256'h9333999993339939DAAAAADDDD22AAA2DDD29DDDAA2DDDDDD222AAA22D922222;
defparam prom_inst_2.INIT_RAM_1B = 256'h933639993E33E9992222AD22D22DDD22ADDDDAA2D22229DA222ADD9DD2D22222;
defparam prom_inst_2.INIT_RAM_1C = 256'h57105434A27911F317250384054054793E4F46E334366034B47FFF46354263E0;
defparam prom_inst_2.INIT_RAM_1D = 256'h843F730F3542EF01543321433C030EEA4AD4FF6FF61FF0EA0934063B2A560013;
defparam prom_inst_2.INIT_RAM_1E = 256'hC3213434113203338F11FFE777043F4028E846904255234C5445763FF76FF524;
defparam prom_inst_2.INIT_RAM_1F = 256'h3FF7539568559565B8A09E45FFF06AAC38092144E8B5F21A9E4208F234548FF8;
defparam prom_inst_2.INIT_RAM_20 = 256'hE2DD92C92EEE0D57A6E6E1C91EA21EFA66E6B2DA019F89FFD3E7E120167DC636;
defparam prom_inst_2.INIT_RAM_21 = 256'h8FE06EAA1BDC5EB58EE7CEC2C2C866E210EE03D5402B06F6ECBDB42816EE1614;
defparam prom_inst_2.INIT_RAM_22 = 256'hCC86DEF8B2B91FEE63C400FEEA7140E5E1652694425716D3EF56C4230315AFA3;
defparam prom_inst_2.INIT_RAM_23 = 256'hEF317163023EEE2F1DEFB923E6E5081AAD54D1D786E26F7190C4C8FF48B509BB;
defparam prom_inst_2.INIT_RAM_24 = 256'hAD0BFFAB0AD00000B0041FAE02F10F00400430E600409B07B060000F000AFD07;
defparam prom_inst_2.INIT_RAM_25 = 256'h20203B801F856062C92005007208004340B070A20DDF0600A30D00D902500010;
defparam prom_inst_2.INIT_RAM_26 = 256'h9107B09D00004D0D009800B908B0000F02C605060A0D90ED6EB001401744B0F8;
defparam prom_inst_2.INIT_RAM_27 = 256'hF7F002FB30A0000382205040006CA0060BEF40100B502A034E00409003C0920A;
defparam prom_inst_2.INIT_RAM_28 = 256'h1CDE5B7233130B8F140E1F5EDD89826AB4A3EFFE52481AA1BD214B05A4CCC78D;
defparam prom_inst_2.INIT_RAM_29 = 256'hFCA15890D83DAE8C20FFC1884B32D49E4C326E4871C5120FB64FF4051E117177;
defparam prom_inst_2.INIT_RAM_2A = 256'hE3442AF09F8016E0C7AC792A4969EC82CD9C1FFC456ABDB4D348F32A9159F692;
defparam prom_inst_2.INIT_RAM_2B = 256'h98D433AC69014868A13F8E2C3ED7182AEF842FEAD5436FF681E93BF9F4512506;
defparam prom_inst_2.INIT_RAM_2C = 256'h166890000CCCCCE7D666666666666664D6666666DDEDA88AA9998433343FA54E;
defparam prom_inst_2.INIT_RAM_2D = 256'hD66666669999DE141989990000BCCCC9E666666666666664E666666FFF0EFE04;
defparam prom_inst_2.INIT_RAM_2E = 256'hB666666666666666C6666CCCC22233251C66990DD000CCE7D666666666666665;
defparam prom_inst_2.INIT_RAM_2F = 256'h5444CCDC78999AAF9666666666666665A666666E1222F0261968880011CCCCC7;
defparam prom_inst_2.INIT_RAM_30 = 256'h23578E88531EEEE5FB29F598654EEEE59E1579A8879ABF4592E940879A93FDDD;
defparam prom_inst_2.INIT_RAM_31 = 256'h4B0311544444AA2E626889ECA96AA4A0A9ACDF10CA9443A395567E862EEC2E75;
defparam prom_inst_2.INIT_RAM_32 = 256'hF07F929BE13578823C6EEE3579BE243FAF36789BBD04AC99F5A44444444BA531;
defparam prom_inst_2.INIT_RAM_33 = 256'h013556A758AABCCD8CD0601454321364C78AE79F2454114BE79DA759CF220031;
defparam prom_inst_2.INIT_RAM_34 = 256'h5FFF00145643344C56AE1311333433395CEF00FF0010B9933762EA2358200000;
defparam prom_inst_2.INIT_RAM_35 = 256'h57C0FCBAAAAA036A7BF1101100C0014A9FF11111100AA46A9CCEF0444451435A;
defparam prom_inst_2.INIT_RAM_36 = 256'h68F716689AAAAAAED91686889989AA9D703566555455095D0F5AAAAAAAA8085C;
defparam prom_inst_2.INIT_RAM_37 = 256'h048CDD187E777777F78C3CBEF010F35D5337B1E36888459E6F164E358AA988AE;
defparam prom_inst_2.INIT_RAM_38 = 256'h7333338808D8880778088830333D33D7088D0003000000877000072822700007;
defparam prom_inst_2.INIT_RAM_39 = 256'h783333D33333388780008888003888027D3388D8333888308000003333333007;
defparam prom_inst_2.INIT_RAM_3A = 256'h80088800888388887880003D300330877033388D83333337200000088830D007;
defparam prom_inst_2.INIT_RAM_3B = 256'h7700077772280000733800883333388720883D33388D03077333330033333337;
defparam prom_inst_2.INIT_RAM_3C = 256'hB344D46434449478D6F8766616737FC666737926D06DFA6633737DA37F5343E3;
defparam prom_inst_2.INIT_RAM_3D = 256'h944443449465444466662907B6B60AA3966F6163756E62636333357773E3333B;
defparam prom_inst_2.INIT_RAM_3E = 256'h4385A44444449F446A63668F6963EA6B66A335BA666056666E337335E7317335;
defparam prom_inst_2.INIT_RAM_3F = 256'h44464346946460547868666386666AE3786666533E666563E53133E03E333A55;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[27:0],dout[15:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 4;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h7777777787677787778777787776776777768887778888777777778688777777;
defparam prom_inst_3.INIT_RAM_01 = 256'h7777776777777777688877778877878876777767777777776888887777777887;
defparam prom_inst_3.INIT_RAM_02 = 256'h6887778877777776777888767887787778777776777777778888888777786887;
defparam prom_inst_3.INIT_RAM_03 = 256'h7777777778867777777788777777777788777677778888877777778877777777;
defparam prom_inst_3.INIT_RAM_04 = 256'h3222533242445523243325364422243453333352433244432524433223332236;
defparam prom_inst_3.INIT_RAM_05 = 256'h3253433022255423333316332324212322552333243124425535345534214444;
defparam prom_inst_3.INIT_RAM_06 = 256'h4322444423764323222234343333322233322235622532344532233346333422;
defparam prom_inst_3.INIT_RAM_07 = 256'h2245544332223543236554333222444452625444222355434222123422233223;
defparam prom_inst_3.INIT_RAM_08 = 256'h3453434453243564352233353335233522453453284332435353323344533445;
defparam prom_inst_3.INIT_RAM_09 = 256'h4433442433445533434355355338333553332332224344233243632433425434;
defparam prom_inst_3.INIT_RAM_0A = 256'h2342344643544334384425524535534343553333322332433233344323434334;
defparam prom_inst_3.INIT_RAM_0B = 256'h2344334438344534443343552323523444532523443433435533333335443423;
defparam prom_inst_3.INIT_RAM_0C = 256'h566A557887577966896658779A5777A677A6688B8A68AA68BA65567AA77AB667;
defparam prom_inst_3.INIT_RAM_0D = 256'h6557658A854457775598876667789587687879B656AAA77A66779A55765555A9;
defparam prom_inst_3.INIT_RAM_0E = 256'h798A66578AA655658AA6577566657855AA6476AA76587876668969AA9A58AAA6;
defparam prom_inst_3.INIT_RAM_0F = 256'h86AA6577A65787586556675557777A8657876787656688AA588A66AA8A759996;
defparam prom_inst_3.INIT_RAM_10 = 256'h5333335595055595559555393330330535509993999999555333359099533335;
defparam prom_inst_3.INIT_RAM_11 = 256'h5533330333333555099955559935659950335505333555330999993333333995;
defparam prom_inst_3.INIT_RAM_12 = 256'h0995559955535550555999303993395559333550533333359999999555390995;
defparam prom_inst_3.INIT_RAM_13 = 256'h5533355559903333533599553333355599553033355093955333339933333335;
defparam prom_inst_3.INIT_RAM_14 = 256'h6666666666666666788888878877778878878777778878887888888788877778;
defparam prom_inst_3.INIT_RAM_15 = 256'h6666666666666666888887777888888877778888788887778888777878877778;
defparam prom_inst_3.INIT_RAM_16 = 256'h6666666666666666788888777788888877787777888777777888888887788888;
defparam prom_inst_3.INIT_RAM_17 = 256'h6665666666666666888887887887778887777888788887788888777778788888;
defparam prom_inst_3.INIT_RAM_18 = 256'h3333333333333333466656635544446646545444445535664666666456644446;
defparam prom_inst_3.INIT_RAM_19 = 256'h3333333333333333666663444666566644445555465553446555344646644446;
defparam prom_inst_3.INIT_RAM_1A = 256'h3333333333333333455555444466555644463444556444444666555664366666;
defparam prom_inst_3.INIT_RAM_1B = 256'h3332333333333333666654664664446654444556466663456665443446466666;
defparam prom_inst_3.INIT_RAM_1C = 256'hEDEEEEEE3213BEFEDDEEBEDDDEDEEEEDEDEDEEDEEEEDDDEEAEEFFFEDDEBEEEDB;
defparam prom_inst_3.INIT_RAM_1D = 256'hDDDFEEBFEDDEDFBEEEEBEEDDDDBEECC3113EFFEFFEEFFE33D3DDDDE3233DBBEE;
defparam prom_inst_3.INIT_RAM_1E = 256'hDDBBDDEEBBBEEEEEEFEEFFDEEEBDDCEBEEDEEDCBDBDDEEEDDDEEEEEDFEEFFDDD;
defparam prom_inst_3.INIT_RAM_1F = 256'hEFFDDDEEEDDD3EEE11DB33DEFFFEE3311143EEEDAEDEDDD333EEEEDEEDDDEFFE;
defparam prom_inst_3.INIT_RAM_20 = 256'h3241431431332223423233143143222142324314324113214333333324314332;
defparam prom_inst_3.INIT_RAM_21 = 256'h3133231424143143313123141324323332314313333433233141432333333323;
defparam prom_inst_3.INIT_RAM_22 = 256'h4143142142433131424325212143323232432413324332433133142323243143;
defparam prom_inst_3.INIT_RAM_23 = 256'h3233133323321332313214341233243114431323323332324223142131433141;
defparam prom_inst_3.INIT_RAM_24 = 256'h9A08A49A08A00000AB09B5A90AA50800505BB04500509B08A050000700059A09;
defparam prom_inst_3.INIT_RAM_25 = 256'h60505BA09A5BA0BA55500600AA05509580505095058408B08908008905A00AA0;
defparam prom_inst_3.INIT_RAM_26 = 256'hA508A09A0000BA0A009500AA0540000509A509050908504859B009909959908B;
defparam prom_inst_3.INIT_RAM_27 = 256'hA58005AA5090000A59B09560008550060AA4905008A09509A40990800BA09B08;
defparam prom_inst_3.INIT_RAM_28 = 256'h89AAA997A9A9A998C999BAA999999CBAAA9A9DAB9998BA9A98DAA9AA999A9AA8;
defparam prom_inst_3.INIT_RAM_29 = 256'hACAA999ABA999A99AAA9CB9999A899A7899989B9AAA9F9A88B89A999BABB9B9A;
defparam prom_inst_3.INIT_RAM_2A = 256'h7999C99A999A9AA999E99ABBA9B8A6AAA9A9B99999A99A989AA998D9AB9AABAA;
defparam prom_inst_3.INIT_RAM_2B = 256'h899AA9B9B8AD89A9A99A97A8A99A99AA9A9AAABAB99978AA99AA99987A9AB9AB;
defparam prom_inst_3.INIT_RAM_2C = 256'hBDDDDEEEEDDDDDDBBEEEEEEEEEEEEEECBEEEEEEEEEEEEEECBBBBBCCCCCCBBBBB;
defparam prom_inst_3.INIT_RAM_2D = 256'hBEEEEEEEEEEEEEFCBDDDDDEEEEDDDDDBBEEEEEEEEEEEEEECBEEEEEEEEEFEEEFC;
defparam prom_inst_3.INIT_RAM_2E = 256'hBEEEEEEEEEEEEEECBEEEEEEEEFFFFFFCBDDDDDEDDEEEDDDBBEEEEEEEEEEEEEEC;
defparam prom_inst_3.INIT_RAM_2F = 256'hBBBBBBBBBBBBBBBBBEEEEEEEEEEEEEECBEEEEEEEFFFFEFFCBDDDDDEEEEDDDDDB;
defparam prom_inst_3.INIT_RAM_30 = 256'h3444445555566664234445555556666434555555555555643544443333332222;
defparam prom_inst_3.INIT_RAM_31 = 256'h3344444444444563344444444444455434444455444445543444445554445654;
defparam prom_inst_3.INIT_RAM_32 = 256'h2444566667777775345555666666777434555555556646642334444444464664;
defparam prom_inst_3.INIT_RAM_33 = 256'h3333333333333333222334555555555423333455666666642333456666777775;
defparam prom_inst_3.INIT_RAM_34 = 256'hBDDDEEEEEEEEEEEBBDDDEEEEEEEEEEEBBDDDEEDDEEEEDDDBBCCCBBBBBBBAAAAA;
defparam prom_inst_3.INIT_RAM_35 = 256'hBDDEDDDDDDDDEEEBBDDEEEEEEEDEEEEBBDDEEEEEEEEDDEEBBDDDDEEEEEEEEEEB;
defparam prom_inst_3.INIT_RAM_36 = 256'hACCDEEEEEEEEEEEBADEEEEEEEEEEEEEBBEEEEEEEEEEEEEEBBCDDDDDDDDDEEEEB;
defparam prom_inst_3.INIT_RAM_37 = 256'hBBBBBBCBBBBBBBBB9BBBCCDDDEEEDEEBACCCCDDEEEEEEEEBABCCDDEEEEEEEEEB;
defparam prom_inst_3.INIT_RAM_38 = 256'h8AAAAAAABA9AAAB88ABAAAABAAA9AA988AA9BBBABBBBBBA88888889799888888;
defparam prom_inst_3.INIT_RAM_39 = 256'h8AAAAA9AAAAAAAA87BBBAAAABBAAAAB989AAAA9AAAAAAAA87BBBBBAAAAAAABB8;
defparam prom_inst_3.INIT_RAM_3A = 256'h7BBAAABBAAAAAAA78AABBBA9ABBAABA88BAAAAA9AAAAAAA89BBBBBBAAAAB9BB8;
defparam prom_inst_3.INIT_RAM_3B = 256'h88888888899788888AAABBAAAAAAAAA89BAAA9AAAAA9BAB88AAAAABBAAAAAAA8;
defparam prom_inst_3.INIT_RAM_3C = 256'h8888988888889888333393333334923333349333233493334444934443449434;
defparam prom_inst_3.INIT_RAM_3D = 256'h9888888898888888933333349323332493323334933234349444444494344443;
defparam prom_inst_3.INIT_RAM_3E = 256'h8888988888889788333493323234933333349333333493333444944444449444;
defparam prom_inst_3.INIT_RAM_3F = 256'h9888888898888888933333349333332493333334923333349444444493444444;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[27:0],dout[19:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 4;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hF44444FFFF8FFFFFFFFFFF4F4448448F4FF8FFF444FFFFFFF4444FF8FFF4444F;
defparam prom_inst_4.INIT_RAM_01 = 256'hFF44448444444FFF8FFFFFFFFF4F0FFFF844FF8F444FFF448FFFFF4444444FFF;
defparam prom_inst_4.INIT_RAM_02 = 256'h8FFFFFFFFFF4FFF8FFFFFF484FF44FFFFF444FF8F444444FFFFFFFFFFF4F8FFF;
defparam prom_inst_4.INIT_RAM_03 = 256'hFF444FFFFFF84444F44FFFFF44444FFFFFFF48444FFFFFFFF44444FF4444444F;
defparam prom_inst_4.INIT_RAM_04 = 256'hC3047D9A05E2067E658095146CF2818F7151D5D39D7C0ACB9630F66F0E67AA8D;
defparam prom_inst_4.INIT_RAM_05 = 256'hF67851268FD55843E1BF6AE731DF9455E6283CA038145865F719F1C76D1D1DAD;
defparam prom_inst_4.INIT_RAM_06 = 256'h99DADDEA71CBC01715DE29E31559E53EEC8CBA86F9C02BC43DF3CAFEA5145742;
defparam prom_inst_4.INIT_RAM_07 = 256'hF01CA9A78E423716163F7EB3F465FFDE6F7551950058737283791772FDAE5DEC;
defparam prom_inst_4.INIT_RAM_08 = 256'h5C55C5CC55DC55CC55DD55555555D555DDC55C55D7C55DC555555D55CC555CC5;
defparam prom_inst_4.INIT_RAM_09 = 256'hCC55CCDC55CC5555C5C55555555755555555D55DDDC5CCD55DC5C5DC55CD5C5C;
defparam prom_inst_4.INIT_RAM_0A = 256'hD5CD5CCCC55CC55C57CCD55DC55555C5C55555555DD55DC55D555CC5D5C5C55C;
defparam prom_inst_4.INIT_RAM_0B = 256'hD5CC55CC575CC55CCC55C555D5D55D5CCC55D5D5CC5855C55555555555CC5CD5;
defparam prom_inst_4.INIT_RAM_0C = 256'h322586FF1F61DB22372465FF292FFA02FF332ED06977C92906DA24E290F9024D;
defparam prom_inst_4.INIT_RAM_0D = 256'h7D323D1796CD6479AE18DF222EA2CE7787FFFEF862D2E2CFF2FFA950F8666699;
defparam prom_inst_4.INIT_RAM_0E = 256'hF15F22132E22A61629910FFA9220F9B2992EFC99260DF7F225CBC0996CD19992;
defparam prom_inst_4.INIT_RAM_0F = 256'h129390FF376F7746566C2FCFDEF4F2C66F8A2D4460187E62A449229BF3D979E2;
defparam prom_inst_4.INIT_RAM_10 = 256'h7333337777777777777777373337337737777773777777777333377777733337;
defparam prom_inst_4.INIT_RAM_11 = 256'h7733337333333777777777777737377777337777333777337777773333333777;
defparam prom_inst_4.INIT_RAM_12 = 256'h7777777777737777777777373773377777333777733333377777777777377777;
defparam prom_inst_4.INIT_RAM_13 = 256'h7733377777773333733777773333377777773733377773777333337733333337;
defparam prom_inst_4.INIT_RAM_14 = 256'h44BBBB4444444BBB9BBB1BB8117777BB9B171777771181BB9BBBBBB71BB7777B;
defparam prom_inst_4.INIT_RAM_15 = 256'h44BBBB444BBBBB44BBBBB8779BBB1BBB777711119B111877B111877B9BB7777B;
defparam prom_inst_4.INIT_RAM_16 = 256'h4BBB44444BBB44B49111117777BB111B977B877711B777779BBB111BB78BBBBB;
defparam prom_inst_4.INIT_RAM_17 = 256'h4BB1B444B8BB8444BBBB17BB9BB777BB1777711B9BBBB871BBB177879B7BBBBB;
defparam prom_inst_4.INIT_RAM_18 = 256'hEE4444EEEEEEE4444888088E00444488480404444400E0884888888408844448;
defparam prom_inst_4.INIT_RAM_19 = 256'hEE4444EEE44444EE88888E44488808884444000048000E448000E44848844448;
defparam prom_inst_4.INIT_RAM_1A = 256'hE444EEEEE444EE4E40000044448800084448E444008444444888000884E88888;
defparam prom_inst_4.INIT_RAM_1B = 256'hE44D4EEE42442EEE88880488488444880444400848888E40888044E448488888;
defparam prom_inst_4.INIT_RAM_1C = 256'h9BCD05A5699C8EFA96BA4C6A6CAAF609A8BFCADE0BF24BBC6D7FFFABDABDEAC4;
defparam prom_inst_4.INIT_RAM_1D = 256'h6D8FFB9F8AC5AF39A7737ABD658B65ADC8BAFFAFFAAFFD1A6C6AD88E9BB144A4;
defparam prom_inst_4.INIT_RAM_1E = 256'hFA29E1BB9969D78A8F38FFAFFF49970B6AF19A9AABAA8A5CEA192DCFFAEFF3C1;
defparam prom_inst_4.INIT_RAM_1F = 256'hFFF6D1DAACCFCBA672D3CAC7FFFAAFC8AE9B44CA3DBB2C8D0E956A9BA3AAAFF9;
defparam prom_inst_4.INIT_RAM_20 = 256'h25C083F831223E889D2D22F821934FBD5D2DA3091482BA02C42822314580B749;
defparam prom_inst_4.INIT_RAM_21 = 256'h9221D2D94A0B61A6912A72F1F3D77D232321F406513A17B72FA0A55927222745;
defparam prom_inst_4.INIT_RAM_22 = 256'hBF770DBBA5AA222156B53FB1FD625328245655C5554829C42267F3543444B294;
defparam prom_inst_4.INIT_RAM_23 = 256'h2042A274334F123B2020E8321D26372DDC4502E89D237B8483D5F7025BA61CAE;
defparam prom_inst_4.INIT_RAM_24 = 256'hAD0BFFAB0AD00000B0041FAE02F10F00400430E600409B07B060000F000AFD07;
defparam prom_inst_4.INIT_RAM_25 = 256'h20203B801F856062C92005007208004340B070A20DDF0600A30D00D902500010;
defparam prom_inst_4.INIT_RAM_26 = 256'h9107B09D00004D0D009800B908B0000F02C605060A0D90ED6EB001401744B0F8;
defparam prom_inst_4.INIT_RAM_27 = 256'hF7F002FB30A0000382205040006CA0060BEF40100B502A034E00409003C0920A;
defparam prom_inst_4.INIT_RAM_28 = 256'h84EFC2FA4A9970E7CC8FCAC65500FE2635236FAFCAC4B5272451507C2C4D578E;
defparam prom_inst_4.INIT_RAM_29 = 256'hAA59C0474EA52A04D7A57C0FC0B85F36C4B8E6A0173CF88724CBAC77C9CCFCFE;
defparam prom_inst_4.INIT_RAM_2A = 256'h3ACCA25705F7DF9740B4F0A6F11093493D548554C722281B53FE5AEC3CC4B139;
defparam prom_inst_4.INIT_RAM_2B = 256'h00543A64118FB0DE59FA0481B6939FD69A0D9A958CCAD7A8E995A05F7AB97C72;
defparam prom_inst_4.INIT_RAM_2C = 256'h166890000CCCCCE7D666666666666664D6666666DDEDA88AA9998433343FA54E;
defparam prom_inst_4.INIT_RAM_2D = 256'hD66666669999DE141989990000BCCCC9E666666666666664E666666FFF0EFE04;
defparam prom_inst_4.INIT_RAM_2E = 256'hB666666666666666C6666CCCC22233251C66990DD000CCE7D666666666666665;
defparam prom_inst_4.INIT_RAM_2F = 256'h5444CCDC78999AAF9666666666666665A666666E1222F0261968880011CCCCC7;
defparam prom_inst_4.INIT_RAM_30 = 256'hF887889BDFDEEEE2E1369A8ABCCEEEE0C33566346775EAA8CDC96279E0C4B1DF;
defparam prom_inst_4.INIT_RAM_31 = 256'hE17BB73111119AD4E38CDBA998599AC3189ABB9999911DE2255678ABCDEBDED1;
defparam prom_inst_4.INIT_RAM_32 = 256'hCE4D7CBCEFEEEDD33F7DEEEFFEDDEEC3E7ADFFEDCBBB9EA389F11111111D9DB4;
defparam prom_inst_4.INIT_RAM_33 = 256'hF37BCD1DD01246784AC0701356877BD5968C0748CEEEBCF5B46C828ACFFDCCE4;
defparam prom_inst_4.INIT_RAM_34 = 256'hF33344589A877885FCF2575577787773F123443344540EEDDFEA74CDF2CDDDDD;
defparam prom_inst_4.INIT_RAM_35 = 256'hFD14310FFFFF47A4103554554414458433355555544FF8A43112348888958794;
defparam prom_inst_4.INIT_RAM_36 = 256'h205D5AABCDDDDDD78E5ABABBCCBCDDC61479AA9998994C96B5BFFFFFFFFB4B95;
defparam prom_inst_4.INIT_RAM_37 = 256'hBE25669217111111C125B302345437961BBF2727ABBB89C7289EA279BDDCBBD7;
defparam prom_inst_4.INIT_RAM_38 = 256'h7333338808D8880778088830333D33D7088D0003000000877000072822700007;
defparam prom_inst_4.INIT_RAM_39 = 256'h783333D33333388780008888003888027D3388D8333888308000003333333007;
defparam prom_inst_4.INIT_RAM_3A = 256'h80088800888388887880003D300330877033388D83333337200000088830D007;
defparam prom_inst_4.INIT_RAM_3B = 256'h7700077772280000733800883333388720883D33388D03077333330033333337;
defparam prom_inst_4.INIT_RAM_3C = 256'h18AA3ACA8AAAFACEE509D555F566DCD55566D9259D525A5566B6DEE6B0769606;
defparam prom_inst_4.INIT_RAM_3D = 256'hFAAAA8AAFAC9AAAAB55529DE1575DC76F55D5F56D35B5556A66668BBD606666C;
defparam prom_inst_4.INIT_RAM_3E = 256'hA8E90AAAAAAAF5AA5A56A59C55563C5C55C683CA555295555366D6683B63D668;
defparam prom_inst_4.INIT_RAM_3F = 256'h9AACA8ACFACAC69AD7595556C5555AB6D75555367B5553564763663270666E87;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[27:0],dout[23:20]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 4;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h7777777787677787778777787776776777768887778888777777778688777777;
defparam prom_inst_5.INIT_RAM_01 = 256'h7777776777777777688877778877878876777767777777776888887777777887;
defparam prom_inst_5.INIT_RAM_02 = 256'h6887778877777776777888767887787778777776777777778888888777786887;
defparam prom_inst_5.INIT_RAM_03 = 256'h7777777778867777777788777777777788777677778888877777778877777777;
defparam prom_inst_5.INIT_RAM_04 = 256'h9999B998B9ABCB999A9A8BACAA898B9ABAAA99B9A998BAA98B9BA9989999889C;
defparam prom_inst_5.INIT_RAM_05 = 256'h99B9BAA7888BBA9A9A998C999A8A889A89BB999A9AA89AA9BBAB9BBBAA97BAAA;
defparam prom_inst_5.INIT_RAM_06 = 256'hA988AAAA9ADCAA999988AA9BAAA999989998889BC88CA89AAB998999ACAAAA99;
defparam prom_inst_5.INIT_RAM_07 = 256'h89BBBAA99899ABB99ACBBA9A9999AAAAB8C9BBAA9999BBAAA998899B8889A889;
defparam prom_inst_5.INIT_RAM_08 = 256'h5685656685365866583355585558355833685685386553658585535566855668;
defparam prom_inst_5.INIT_RAM_09 = 256'h6655663655668855656588588558555885553553336566355365653655638656;
defparam prom_inst_5.INIT_RAM_0A = 256'h3563566665866556586638836858856565885555533553655355566535656556;
defparam prom_inst_5.INIT_RAM_0B = 256'h3566556658566856665565883535835666853835665555658855555558665635;
defparam prom_inst_5.INIT_RAM_0C = 256'h566A557887577966896658779A5777A677A6688B8A68AA68BA65567AA77AB667;
defparam prom_inst_5.INIT_RAM_0D = 256'h6557658A854457775598876667789587687879B656AAA77A66779A55765555A9;
defparam prom_inst_5.INIT_RAM_0E = 256'h798A66578AA655658AA6577566657855AA6476AA76587876668969AA9A58AAA6;
defparam prom_inst_5.INIT_RAM_0F = 256'h86AA6577A65787586556675557777A8657876787656688AA588A66AA8A759996;
defparam prom_inst_5.INIT_RAM_10 = 256'h5333335595055595559555393330330535509993999999555333359099533335;
defparam prom_inst_5.INIT_RAM_11 = 256'h5533330333333555099955559935659950335505333555330999993333333995;
defparam prom_inst_5.INIT_RAM_12 = 256'h0995559955535550555999303993395559333550533333359999999555390995;
defparam prom_inst_5.INIT_RAM_13 = 256'h5533355559903333533599553333355599553033355093955333339933333335;
defparam prom_inst_5.INIT_RAM_14 = 256'h9988889999999888ACCCCCCACCBBBBCCACCBCBBBBBCCACCCACCCCCCBCCCBBBBC;
defparam prom_inst_5.INIT_RAM_15 = 256'h9988889998888899CCCCCABBACCCCCCCBBBBCCCCACCCCABBCCCCABBCACCBBBBC;
defparam prom_inst_5.INIT_RAM_16 = 256'h9888999998889989ACCCCCBBBBCCCCCCABBCABBBCCCBBBBBACCCCCCCCBACCCCC;
defparam prom_inst_5.INIT_RAM_17 = 256'h9888899989889999CCCCCBCCACCBBBCCCBBBBCCCACCCCABCCCCCBBABACBCCCCC;
defparam prom_inst_5.INIT_RAM_18 = 256'h5555555555555555899999959988889989989888889959998999999899988889;
defparam prom_inst_5.INIT_RAM_19 = 256'h5555555555555555999995888999999988889999899995889999588989988889;
defparam prom_inst_5.INIT_RAM_1A = 256'h5555555555555555899999888899999988895888999888888999999998599999;
defparam prom_inst_5.INIT_RAM_1B = 256'h5553555556556555999998998998889998888999899995899999885889899999;
defparam prom_inst_5.INIT_RAM_1C = 256'hEDEEFEEE3113BEFEDDEEBEDDDEDEEEFDEEEEEEEEEEEDDDEEBEEFFFEDDEBEEEEB;
defparam prom_inst_5.INIT_RAM_1D = 256'hDDDFEEBFEDDEEFBEEEEBEEDDDEBEEDD3113EFFEFFEEFFE43D3DDDDE3133EBBEE;
defparam prom_inst_5.INIT_RAM_1E = 256'hDDBBDEEEBBBEEEEEEFEEFFEEEEBDDDFBEEEFEDDBDBDDEEEEDDFEEEEDFEEFFDDD;
defparam prom_inst_5.INIT_RAM_1F = 256'hEFFDDDEEEDDD3EEE12DB33DEFFFEE3311133EEEDBEEEFDD343EEEEEEEEDDEFFE;
defparam prom_inst_5.INIT_RAM_20 = 256'h6373752753663435736365275375344273637537537325537565655537537553;
defparam prom_inst_5.INIT_RAM_21 = 256'h5365362737375375536246272547536553636535555755456273753555665535;
defparam prom_inst_5.INIT_RAM_22 = 256'h7275374273755363737537434275536363753725537553756355273535375375;
defparam prom_inst_5.INIT_RAM_23 = 256'h6555255535543654536527573365375227753545536554537345275352755272;
defparam prom_inst_5.INIT_RAM_24 = 256'h9A08A49A08A00000AB09B5A90AA50800505BB04500509B08A050000700059A09;
defparam prom_inst_5.INIT_RAM_25 = 256'h60505BA09A5BA0BA55500600AA05509580505095058408B08908008905A00AA0;
defparam prom_inst_5.INIT_RAM_26 = 256'hA508A09A0000BA0A009500AA0540000509A509050908504859B009909959908B;
defparam prom_inst_5.INIT_RAM_27 = 256'hA58005AA5090000A59B09560008550060AA4905008A09509A40990800BA09B08;
defparam prom_inst_5.INIT_RAM_28 = 256'hBDDDDDCADCDCDDCCECCCDDDDDDDDCEEDEDDDDFDDCCCBDDDDDCFDDDDDDCDDDDDB;
defparam prom_inst_5.INIT_RAM_29 = 256'hDEDDCDCDFDCDDDDDCDDDFDDCCDDBDBDBBDCCBDEDDDECFCDCCEBCDCCCDDDDCDCD;
defparam prom_inst_5.INIT_RAM_2A = 256'hBCCCFDDDDDCDBDDCDDFDCEEECDECDADDECDDEDDDCCDDDDDBDDCCDBFCDDCDDEDD;
defparam prom_inst_5.INIT_RAM_2B = 256'hCDDDDCEDECDFBDDCDCBDDBDCDDCDCCCDCDDDDDEDECCCACDDCCDDCDDBBDCDECDE;
defparam prom_inst_5.INIT_RAM_2C = 256'hBDDDDEEEEDDDDDDBBEEEEEEEEEEEEEECBEEEEEEEEEEEEEECBBBBBCCCCCCBBBBB;
defparam prom_inst_5.INIT_RAM_2D = 256'hBEEEEEEEEEEEEEFCBDDDDDEEEEDDDDDBBEEEEEEEEEEEEEECBEEEEEEEEEFEEEFC;
defparam prom_inst_5.INIT_RAM_2E = 256'hBEEEEEEEEEEEEEECBEEEEEEEEFFFFFFCBDDDDDEDDEEEDDDBBEEEEEEEEEEEEEEC;
defparam prom_inst_5.INIT_RAM_2F = 256'hBBBBBBBBBBBBBBBBBEEEEEEEEEEEEEECBEEEEEEEFFFFEFFCBDDDDDEEEEDDDDDB;
defparam prom_inst_5.INIT_RAM_30 = 256'hCFFFFFFFFFFFFFFDCFFFFFFFFFFFFFFDCFFFFFFFFFFFEEECCDDDDDCCCDCCBBAA;
defparam prom_inst_5.INIT_RAM_31 = 256'hCFFFFFFFFFFFFFFDCFFFFFFFFFFFFFFDDFFFFFFFFFFFFFFDDFFFFFFFFFFFFFFD;
defparam prom_inst_5.INIT_RAM_32 = 256'hBDEEFFFFFFFFFFFDCEFFFFFFFFFFFFFDCFFFFFFFFFFFFFFDCEEFFFFFFFFFFFFD;
defparam prom_inst_5.INIT_RAM_33 = 256'hBCCCCCDCCDDDDDDDBCCDDEFFFFFFFFFDBDDDEEFFFFFFFFFDBDDDEFFFFFFFFFFD;
defparam prom_inst_5.INIT_RAM_34 = 256'hBEEEEEEEEEEEEEECBDDEEEEEEEEEEEECBEEEEEEEEEEEEDDBBCCCCCBBBCBAAAAA;
defparam prom_inst_5.INIT_RAM_35 = 256'hBDEEEEEDDDDDEEECCEEEEEEEEEEEEEECCEEEEEEEEEEDDEECCEEEEEEEEEEEEEEC;
defparam prom_inst_5.INIT_RAM_36 = 256'hBDDDEEEEEEEEEEECBDEEEEEEEEEEEEECCEEEEEEEEEEEEEECBDDDDDDDDDDEEEEC;
defparam prom_inst_5.INIT_RAM_37 = 256'hBBCCCCCCCCCCCCCCACCCCDEEEEEEEEECBCCCDDEEEEEEEEECBCCCDEEEEEEEEEEC;
defparam prom_inst_5.INIT_RAM_38 = 256'h8AAAAAAABA9AAAB88ABAAAABAAA9AA988AA9BBBABBBBBBA88888889799888888;
defparam prom_inst_5.INIT_RAM_39 = 256'h8AAAAA9AAAAAAAA87BBBAAAABBAAAAB989AAAA9AAAAAAAA87BBBBBAAAAAAABB8;
defparam prom_inst_5.INIT_RAM_3A = 256'h7BBAAABBAAAAAAA78AABBBA9ABBAABA88BAAAAA9AAAAAAA89BBBBBBAAAAB9BB8;
defparam prom_inst_5.INIT_RAM_3B = 256'h88888888899788888AAABBAAAAAAAAA89BAAA9AAAAA9BAB88AAAAABBAAAAAAA8;
defparam prom_inst_5.INIT_RAM_3C = 256'h9888A888888898884454944434459344444594443346A4445555945555559555;
defparam prom_inst_5.INIT_RAM_3D = 256'h988888889888888894444435A434343594434345944345459555555595555554;
defparam prom_inst_5.INIT_RAM_3E = 256'h8888A88888889888444594434345A44444459444444594444655955565559555;
defparam prom_inst_5.INIT_RAM_3F = 256'h988888889888888894444445944444359444444593444445A555556595555555;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[27:0],dout[27:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 4;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hF44444FFFF8FFFFFFFFFFF4F4448448F4FF8FFF444FFFFFFF4444FF8FFF4444F;
defparam prom_inst_6.INIT_RAM_01 = 256'hFF44448444444FFF8FFFFFFFFF4F0FFFF844FF8F444FFF448FFFFF4444444FFF;
defparam prom_inst_6.INIT_RAM_02 = 256'h8FFFFFFFFFF4FFF8FFFFFF484FF44FFFFF444FF8F444444FFFFFFFFFFF4F8FFF;
defparam prom_inst_6.INIT_RAM_03 = 256'hFF444FFFFFF84444F44FFFFF44444FFFFFFF48444FFFFFFFF44444FF4444444F;
defparam prom_inst_6.INIT_RAM_04 = 256'hE63A38229708C6B281A3C4AFEB78BCEE3782C1BE90CF96CBE5CEB1BF41BADBCE;
defparam prom_inst_6.INIT_RAM_05 = 256'hA9AB8269C4011B74F2F2996A6406C7A636436A536925A4C6A3F8D3728922DB6E;
defparam prom_inst_6.INIT_RAM_06 = 256'hCCEDB9FE8474F34A6A04B22DA4B07A83F89FECB2D1FC5E2029E6FD21A4648C7B;
defparam prom_inst_6.INIT_RAM_07 = 256'h1F0CA87AB48310FC992D5AF407CBAF0143053F25338B31D51688ABA240D2A232;
defparam prom_inst_6.INIT_RAM_08 = 256'h96996966999699C6999999999999999999699699976999699999999966999669;
defparam prom_inst_6.INIT_RAM_09 = 256'h6699669699669999696999999997999999999999996966999969C99699699696;
defparam prom_inst_6.INIT_RAM_0A = 256'h9969966C69966996976699996999996969999999999999699999966999696996;
defparam prom_inst_6.INIT_RAM_0B = 256'h9966996697966996669969999999999666999999669499699999999999669699;
defparam prom_inst_6.INIT_RAM_0C = 256'h322586FF1F61DB22372465FF292FFA02FF332ED06977C92906DA24E290F9024D;
defparam prom_inst_6.INIT_RAM_0D = 256'h7D323D1796CD6479AE18DF222EA2CE7787FFFEF862D2E2CFF2FFA950F8666699;
defparam prom_inst_6.INIT_RAM_0E = 256'hF15F22132E22A61629910FFA9220F9B2992EFC99260DF7F225CBC0996CD19992;
defparam prom_inst_6.INIT_RAM_0F = 256'h129390FF376F7746566C2FCFDEF4F2C66F8A2D4460187E62A449229BF3D979E2;
defparam prom_inst_6.INIT_RAM_10 = 256'h7333337777777777777777373337337737777773777777777333377777733337;
defparam prom_inst_6.INIT_RAM_11 = 256'h7733337333333777777777777737377777337777333777337777773333333777;
defparam prom_inst_6.INIT_RAM_12 = 256'h7777777777737777777777373773377777333777733333377777777777377777;
defparam prom_inst_6.INIT_RAM_13 = 256'h7733377777773333733777773333377777773733377773777333337733333337;
defparam prom_inst_6.INIT_RAM_14 = 256'h55EEEE5555555EEEA777777877888877A778788888778777A777777877788887;
defparam prom_inst_6.INIT_RAM_15 = 256'h55EEEE555EEEEE5577777888A777777788887777A777788877778887A7788887;
defparam prom_inst_6.INIT_RAM_16 = 256'h5EEE55555EEE55E5A777778888777777A887888877788888A777777778877777;
defparam prom_inst_6.INIT_RAM_17 = 256'h5EEEE555EEEEE55577777877A778887778888777A777788777778888A7877777;
defparam prom_inst_6.INIT_RAM_18 = 256'h3399993333333999FCCC4CC344FFFFCCFC4F4FFFFF4434CCFCCCCCCF4CCFFFFC;
defparam prom_inst_6.INIT_RAM_19 = 256'h3399993339999933CCCCC3FFFCCC4CCCFFFF4444FC4443FFC4443FFCFCCFFFFC;
defparam prom_inst_6.INIT_RAM_1A = 256'h3999333339993393F44444FFFFCC444CFFFC3FFF44CFFFFFFCCC444CCF3CCCCC;
defparam prom_inst_6.INIT_RAM_1B = 256'h399C93339C99C333CCCC4FCCFCCFFFCC4FFFF44CFCCCC3F4CCC4FF3FFCFCCCCC;
defparam prom_inst_6.INIT_RAM_1C = 256'hAAD8EA1DC05113FEB95867ACDB2BD78681CAB787A66CB9721B9FFF40BD8CEBA2;
defparam prom_inst_6.INIT_RAM_1D = 256'h79DFA6FF6EBACFA7B9F4AF92BAB81A0DADCDFFBFFA0FFD1AA20B595E0DED66BA;
defparam prom_inst_6.INIT_RAM_1E = 256'h9D40D5DD00C936B9AF4AFFCCCC6FBAC79099C696F1EE293CD2C3D0AAF18FFEAC;
defparam prom_inst_6.INIT_RAM_1F = 256'h4FFC07DAD2A9BAB8CDAACABDFFF9A6F9BFE08B9856AEC7BA2E9AB87AA7B7CFF3;
defparam prom_inst_6.INIT_RAM_20 = 256'hC2CD88C88ECC035D9CCCC7C87E9814EA5CCCA8D9618F8F5FC9CDC78615DDBC96;
defparam prom_inst_6.INIT_RAM_21 = 256'hEFC6CCA91ADBBEABEEC79CC1C827CCC870CEF9DBA68A6CECCCADAA2E7CCC7C1A;
defparam prom_inst_6.INIT_RAM_22 = 256'hBC7CDDE8A2AF7FCE53BA0FEE4A67A0C5C15B259AA24D76C9CFBCC32909140F99;
defparam prom_inst_6.INIT_RAM_23 = 256'hC59777C90894EC8E7DC5B882ECCB077AAC4AD73DECC8CED1802AC75FA8AB69AB;
defparam prom_inst_6.INIT_RAM_24 = 256'hAD0BFFAB0AD00000B0041FAE02F10F00400430E600409B07B060000F000AFD07;
defparam prom_inst_6.INIT_RAM_25 = 256'h20203B801F856062C92005007208004340B070A20DDF0600A30D00D902500010;
defparam prom_inst_6.INIT_RAM_26 = 256'h9107B09D00004D0D009800B908B0000F02C605060A0D90ED6EB001401744B0F8;
defparam prom_inst_6.INIT_RAM_27 = 256'hF7F002FB30A0000382205040006CA0060BEF40100B502A034E00409003C0920A;
defparam prom_inst_6.INIT_RAM_28 = 256'hFA782960D1F0D86C82F9862CBB6869E29F8ECF62302F708E9A7CF8D282A6B127;
defparam prom_inst_6.INIT_RAM_29 = 256'h6E0F360DB51B866A9D6CF866282FBBFC2A1F5C16DE93FFFD9E2762D086886864;
defparam prom_inst_6.INIT_RAM_2A = 256'hB122F8CD8C6D955EA6BA6611B7D7590FA70AECCA20D89481BDB6C1F5F8307DF0;
defparam prom_inst_6.INIT_RAM_2B = 256'h66BFE11AD7FF16360FB66BF81C5EF7825663F66043213C6E605018C7E22FF3DE;
defparam prom_inst_6.INIT_RAM_2C = 256'h166890000CCCCCE7D666666666666664D6666666DDEDA88AA9998433343FA54E;
defparam prom_inst_6.INIT_RAM_2D = 256'hD66666669999DE141989990000BCCCC9E666666666666664E666666FFF0EFE04;
defparam prom_inst_6.INIT_RAM_2E = 256'hB666666666666666C6666CCCC22233251C66990DD000CCE7D666666666666665;
defparam prom_inst_6.INIT_RAM_2F = 256'h5444CCDC78999AAF9666666666666665A666666E1222F0261968880011CCCCC7;
defparam prom_inst_6.INIT_RAM_30 = 256'h9FFFFECDEEDFFFFAAABEFECBBBCFFFF8AFFFFFFEEEEEFED7A0FDABCBAA830A88;
defparam prom_inst_6.INIT_RAM_31 = 256'h9CDDBAEFFFFFFDD8AEDC99FFFFDFFAB7ACCDDDEFFFFFFDEAADDDEEFFFFFDDFFA;
defparam prom_inst_6.INIT_RAM_32 = 256'h689CFFEEFFFFFFFA8EFFFEDDEEFFFFFAAFFEECDDEEEFFFFA87BFFFFFFFFFFFFA;
defparam prom_inst_6.INIT_RAM_33 = 256'hABDFFD2FE0DDEEEE6656CCEFFFFEDDFA9CAACBCDFFFEBBEA8646EFDDFFFFDEFA;
defparam prom_inst_6.INIT_RAM_34 = 256'h0DDD22716B1CC1100A987C77CCC1CCC0038D22DD2272E4400E9A000000000000;
defparam prom_inst_6.INIT_RAM_35 = 256'h0F32D3E999992CB00ED77277223227100DD77777722991B00338D21111671C60;
defparam prom_inst_6.INIT_RAM_36 = 256'h03CF7BB05AAAAAA0047B0B005505AA5002C6BB66616625600C59999999902060;
defparam prom_inst_6.INIT_RAM_37 = 256'h00000050000000000000F2E8D272DC600FFED68CB0001650005908C60AA500A0;
defparam prom_inst_6.INIT_RAM_38 = 256'h7333338808D8880778088830333D33D7088D0003000000877000072822700007;
defparam prom_inst_6.INIT_RAM_39 = 256'h783333D33333388780008888003888027D3388D8333888308000003333333007;
defparam prom_inst_6.INIT_RAM_3A = 256'h80088800888388887880003D300330877033388D83333337200000088830D007;
defparam prom_inst_6.INIT_RAM_3B = 256'h7700077772280000733800883333388720883D33388D03077333330033333337;
defparam prom_inst_6.INIT_RAM_3C = 256'h3BEE5E0EBEEE1CF0DCF2FCCC3CFBFBCCECFBF36C7EC176CCBB5BFDAB5FDBCB2B;
defparam prom_inst_6.INIT_RAM_3D = 256'h1EEEEBEE1E0DCEEEECCC63E75C5CE82B1CCDC3CBF9CACACBEBBBBF55FB2BBBB9;
defparam prom_inst_6.INIT_RAM_3E = 256'hEB0D2CEEEEEE19EEC6CBEC2BCFCB68C9CC8BB996CCC4DCCCE2BBFBBF23B7FBBF;
defparam prom_inst_6.INIT_RAM_3F = 256'hCEE0EBE01EEEE8DEF0C2CCCB0CCCC6ABF0ECCC9BBACCC9CB8DB7BB24B2BBBAFD;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[27:0],dout[31:28]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 4;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h7777777787677787778777787776776777768887778888777777778688777777;
defparam prom_inst_7.INIT_RAM_01 = 256'h7777776777777777688877778877878876777767777777776888887777777887;
defparam prom_inst_7.INIT_RAM_02 = 256'h6887778877777776777888767887787778777776777777778888888777786887;
defparam prom_inst_7.INIT_RAM_03 = 256'h7777777778867777777788777777777788777677778888877777778877777777;
defparam prom_inst_7.INIT_RAM_04 = 256'h5555866575778856575648686755475786665685665477654857765456554459;
defparam prom_inst_7.INIT_RAM_05 = 256'h6575766345588656565649655657445655885666566457658868688867547776;
defparam prom_inst_7.INIT_RAM_06 = 256'h6544776656A96655555567676666655556544458954864677855456679666655;
defparam prom_inst_7.INIT_RAM_07 = 256'h5488877555556875569887566555777785958777555588667554455855466556;
defparam prom_inst_7.INIT_RAM_08 = 256'h79B79799B7597B697B55777B777B577B559B79B758977597B7B7757799B7799B;
defparam prom_inst_7.INIT_RAM_09 = 256'h997799597799BB779797BB7BB778777BB777577555979957759767597795B979;
defparam prom_inst_7.INIT_RAM_0A = 256'h5795799697B9977978995BB59B7BB79797BB7777755775977577799757979779;
defparam prom_inst_7.INIT_RAM_0B = 256'h5799779978799B79997797BB5757B57999B75B5799777797BB7777777B997957;
defparam prom_inst_7.INIT_RAM_0C = 256'h566A557887577966896658779A5777A677A6688B8A68AA68BA65567AA77AB667;
defparam prom_inst_7.INIT_RAM_0D = 256'h6557658A854457775598876667789587687879B656AAA77A66779A55765555A9;
defparam prom_inst_7.INIT_RAM_0E = 256'h798A66578AA655658AA6577566657855AA6476AA76587876668969AA9A58AAA6;
defparam prom_inst_7.INIT_RAM_0F = 256'h86AA6577A65787586556675557777A8657876787656688AA588A66AA8A759996;
defparam prom_inst_7.INIT_RAM_10 = 256'h5333335595055595559555393330330535509993999999555333359099533335;
defparam prom_inst_7.INIT_RAM_11 = 256'h5533330333333555099955559935659950335505333555330999993333333995;
defparam prom_inst_7.INIT_RAM_12 = 256'h0995559955535550555999303993395559333550533333359999999555390995;
defparam prom_inst_7.INIT_RAM_13 = 256'h5533355559903333533599553333355599553033355093955333339933333335;
defparam prom_inst_7.INIT_RAM_14 = 256'hAA9999AAAAAAA999BDDDDDDBDDCCCCDDBDDCDCCCCCDDBDDDBDDDDDDCDDDCCCCD;
defparam prom_inst_7.INIT_RAM_15 = 256'hAA9999AAA99999AADDDDDBCCBDDDDDDDCCCCDDDDBDDDDBCCDDDDBCCDBDDCCCCD;
defparam prom_inst_7.INIT_RAM_16 = 256'hA999AAAAA999AA9ABDDDDDCCCCDDDDDDBCCDBCCCDDDCCCCCBDDDDDDDDCBDDDDD;
defparam prom_inst_7.INIT_RAM_17 = 256'hA9989AAA9A99AAAADDDDDCDDBDDCCCDDDCCCCDDDBDDDDBCDDDDDCCBCBDCDDDDD;
defparam prom_inst_7.INIT_RAM_18 = 256'h77666677777776669BBBBBB7BB9999BB9BB9B99999BB7BBB9BBBBBB9BBB9999B;
defparam prom_inst_7.INIT_RAM_19 = 256'h7766667776666677BBBBB7999BBBBBBB9999BBBB9BBBB799BBBB799B9BB9999B;
defparam prom_inst_7.INIT_RAM_1A = 256'h76667777766677679BBBBB9999BBBBBB999B7999BBB999999BBBBBBBB97BBBBB;
defparam prom_inst_7.INIT_RAM_1B = 256'h7664677767667777BBBBB9BB9BB999BBB9999BBB9BBBB79BBBBB99799B9BBBBB;
defparam prom_inst_7.INIT_RAM_1C = 256'hEDEEEEFE3214BEFEDDEEBEDDDEEEEEEDEFEEEEEEEEEDDDEFBEEFFFEEDEBEEEEB;
defparam prom_inst_7.INIT_RAM_1D = 256'hDDDFEEBFEDDEEFBEEEEBEEDDDEBEEDE3113EFFEFFEFFFE43D4EDDDE3233DBBEE;
defparam prom_inst_7.INIT_RAM_1E = 256'hDDBBDDEEBBBEEEEEEFEEFFEEEEBDDDEBEFEEEDDBDBDDEEEEDDEEEFEEFFEFFDDD;
defparam prom_inst_7.INIT_RAM_1F = 256'hFFFDEDEEEEDD3EEE11DB33DEFFFEE3311134EEEDBEEEEDD343EEEEEEEDDDEFFE;
defparam prom_inst_7.INIT_RAM_20 = 256'h7493963963774646947476396396465394749639649336639676766649639664;
defparam prom_inst_7.INIT_RAM_21 = 256'h6376473949396396637357393669647664738636666966567393964666776646;
defparam prom_inst_7.INIT_RAM_22 = 256'h9396395394966373949649536396647474964936649664967366394646497396;
defparam prom_inst_7.INIT_RAM_23 = 256'h7666366646663765637639693476496339963666647665649466396363966393;
defparam prom_inst_7.INIT_RAM_24 = 256'h9A08A49A08A00000AB09B5A90AA50800505BB04500509B08A050000700059A09;
defparam prom_inst_7.INIT_RAM_25 = 256'h60505BA09A5BA0BA55500600AA05509580505095058408B08908008905A00AA0;
defparam prom_inst_7.INIT_RAM_26 = 256'hA508A09A0000BA0A009500AA0540000509A509050908504859B009909959908B;
defparam prom_inst_7.INIT_RAM_27 = 256'hA58005AA5090000A59B09560008550060AA4905008A09509A40990800BA09B08;
defparam prom_inst_7.INIT_RAM_28 = 256'hBDEEEDDBDDDDDDDCFDCDEEEDDDDDDFEEEDDDDFEEDDDBEEDDDCFDDDDEDDDEDEEC;
defparam prom_inst_7.INIT_RAM_29 = 256'hEEEDDDDDFEDDDEDDDDEDFEDDDDEBDCDBCDDCCDFDDDEDFCDCCECDEDCDEEEEDEDE;
defparam prom_inst_7.INIT_RAM_2A = 256'hBDDDFDDDDDDDCEECDDFDDEFFDDECEAEDEDEDEDDDDDDDDEDCDDDDDCFDDEDEEEDE;
defparam prom_inst_7.INIT_RAM_2B = 256'hCDDDDDFDECDFCDEDECCEDBDCEDDDCDDEDEDEDEFEFDDDBCEDDDEEDDDCBEDDEDDE;
defparam prom_inst_7.INIT_RAM_2C = 256'hBDDDDEEEEDDDDDDBBEEEEEEEEEEEEEECBEEEEEEEEEEEEEECBBBBBCCCCCCBBBBB;
defparam prom_inst_7.INIT_RAM_2D = 256'hBEEEEEEEEEEEEEFCBDDDDDEEEEDDDDDBBEEEEEEEEEEEEEECBEEEEEEEEEFEEEFC;
defparam prom_inst_7.INIT_RAM_2E = 256'hBEEEEEEEEEEEEEECBEEEEEEEEFFFFFFCBDDDDDEDDEEEDDDBBEEEEEEEEEEEEEEC;
defparam prom_inst_7.INIT_RAM_2F = 256'hBBBBBBBBBBBBBBBBBEEEEEEEEEEEEEECBEEEEEEEFFFFEFFCBDDDDDEEEEDDDDDB;
defparam prom_inst_7.INIT_RAM_30 = 256'hEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFEEEEEEEEEEEDDD;
defparam prom_inst_7.INIT_RAM_31 = 256'hEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFE;
defparam prom_inst_7.INIT_RAM_32 = 256'hEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFE;
defparam prom_inst_7.INIT_RAM_33 = 256'hFFFFFFFEEFEEEEEEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFE;
defparam prom_inst_7.INIT_RAM_34 = 256'h0777888999988990056788888889888007778877888866600110000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0578776666668890067888888878889007788888888669900777789999989890;
defparam prom_inst_7.INIT_RAM_36 = 256'h0235899AAAAAAAA00689A9AAAAAAAAA00889999999998A9003566666666A8A90;
defparam prom_inst_7.INIT_RAM_37 = 256'h00000000000000000000036778887890000124789AAA99A000015789AAAAAAA0;
defparam prom_inst_7.INIT_RAM_38 = 256'h8AAAAAAABA9AAAB88ABAAAABAAA9AA988AA9BBBABBBBBBA88888889799888888;
defparam prom_inst_7.INIT_RAM_39 = 256'h8AAAAA9AAAAAAAA87BBBAAAABBAAAAB989AAAA9AAAAAAAA87BBBBBAAAAAAABB8;
defparam prom_inst_7.INIT_RAM_3A = 256'h7BBAAABBAAAAAAA78AABBBA9ABBAABA88BAAAAA9AAAAAAA89BBBBBBAAAAB9BB8;
defparam prom_inst_7.INIT_RAM_3B = 256'h88888888899788888AAABBAAAAAAAAA89BAAA9AAAAA9BAB88AAAAABBAAAAAAA8;
defparam prom_inst_7.INIT_RAM_3C = 256'hA999B9A99999B99A8788A7777779A6877779A877667BB87799A9A8A9A899A999;
defparam prom_inst_7.INIT_RAM_3D = 256'hB9999999B9A99999A777786AB7676869B7767779A7767979A99999AAA9999998;
defparam prom_inst_7.INIT_RAM_3E = 256'h99A9B9999999B9997879A7867579B8787789A7887779A7777B99A999BA99A999;
defparam prom_inst_7.INIT_RAM_3F = 256'hA99A999AB9999999A8787779B7777869A8777779A6777779B99999B9A9999A99;

endmodule //texture_rom
