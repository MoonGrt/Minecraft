//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Tue Sep 23 22:52:19 2025

module map_ram (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [3:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [14:0] ada;
input [3:0] din;
input [14:0] adb;

wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [1:1] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [1:1] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [2:2] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [2:2] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [3:3] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [3:3] sdpb_inst_7_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0000010100000101000001010000010100000101000003010000010100000101;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h0000010100000101000001010000010100000101000001010000030100000101;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h0000010100000101000001010000010100000101000001010000010100000101;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h0000010100000101000001010000010100000101000001010000010100003F01;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h0000010100000101000001010000010100000101000001010000010100000101;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h0000010100000101000001010000010100000101000001010000010100000101;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_0B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_0D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_17 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_19 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_22 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_23 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_24 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_25 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_26 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_27 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h0000017E0000017E0000017E0000017E0000017E0000037E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_2A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_2E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_2F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_32 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_35 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_37 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_3C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_3D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_02 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E00003F7E;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_05 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_06 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_07 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_09 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_0A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_0B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_0C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_0E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_11 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_13 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_14 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h0000017E0000017E0000017E0000037E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_18 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_19 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_1A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_1B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_1C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_1D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_1E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_1F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_20 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_23 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_24 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_26 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_2E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_30 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_31 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_32 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_33 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_38 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_3A = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;
defparam sdpb_inst_3.INIT_RAM_3F = 256'h0000017E0000017E0000017E0000017E0000017E0000017E0000017E0000017E;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000020000000000;
defparam sdpb_inst_4.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000003E00;
defparam sdpb_inst_5.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_12 = 256'h0000000000000000000000000000020000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_16 = 256'h0000000000000000000000000000020000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000002000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000020000000000;
defparam sdpb_inst_6.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_39 = 256'h0000200000002000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000020000000200000002000;
defparam sdpb_inst_6.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3D = 256'h0000E00000002000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000020000000E0000000E000;
defparam sdpb_inst_6.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_01 = 256'h0000E00000002000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000020000000E0000000C000;
defparam sdpb_inst_7.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_05 = 256'h0000E00000002000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000020000000E0000000E000;
defparam sdpb_inst_7.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_09 = 256'h0000200000002000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000020000000200000002000;
defparam sdpb_inst_7.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_12 = 256'h0000000000000000000000000000020000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_16 = 256'h0000000000000000000000000000020000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(sdpb_inst_2_dout[1]),
  .I1(sdpb_inst_3_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(sdpb_inst_4_dout[2]),
  .I1(sdpb_inst_5_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(sdpb_inst_6_dout[3]),
  .I1(sdpb_inst_7_dout[3]),
  .S0(dff_q_0)
);
endmodule //map_ram
